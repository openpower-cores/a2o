// © IBM Corp. 2020
// This softcore is licensed under and subject to the terms of the CC-BY 4.0
// license (https://creativecommons.org/licenses/by/4.0/legalcode). 
// Additional rights, including the right to physically implement a softcore 
// that is compliant with the required sections of the Power ISA 
// Specification, will be available at no cost via the OpenPOWER Foundation. 
// This README will be updated with additional information when OpenPOWER's 
// license is available.

`timescale 1 ns / 1 ns

//-------------------------------------------------------------------

//-------------------------------------------------------------------

`include "tri_a2o.vh"

module iuq_axu_fu_dec(
   input [0:`NCLK_WIDTH-1]   nclk,
   //-------------------------------------------------------------------
   inout                     vdd,
   inout                     gnd,
   //-------------------------------------------------------------------

   input                     i_dec_si,
   output                    i_dec_so,

   input                     pc_iu_sg_2,
   input                     pc_iu_func_sl_thold_2,
   input                     clkoff_b,
   input                     act_dis,
   input                     tc_ac_ccflush_dc,
   input                     d_mode,
   input                     delay_lclkr,
   input                     mpw1_b,
   input                     mpw2_b,

   input                     iu_au_iu4_isram,

   // AXU interface signals---------------------------------------------
   input                     iu_au_iu4_instr_v,
   input [0:31]              iu_au_iu4_instr,
   input [0:3]               iu_au_iu4_ucode_ext,		// TABC
   input [0:2]               iu_au_iu4_ucode,
   input                     iu_au_iu4_2ucode,
   input                     iu_au_ucode_restart,

   input [0:7]               iu_au_config_iucr,		// 0: graphics mode, 1: disable axu bypass

   // out to AXU
   output                    au_iu_iu4_i_dec_b,		// decoded a valid FU instruction (inverted) 0509
   output [0:2]              au_iu_iu4_ucode,

   output                    au_iu_iu4_t1_v,
   output [0:2]              au_iu_iu4_t1_t,
   output [0:`GPR_POOL_ENC-1] au_iu_iu4_t1_a,

   output                    au_iu_iu4_t2_v,
   output [0:`GPR_POOL_ENC-1] au_iu_iu4_t2_a,
   output [0:2]              au_iu_iu4_t2_t,

   output                    au_iu_iu4_t3_v,
   output [0:`GPR_POOL_ENC-1] au_iu_iu4_t3_a,
   output [0:2]              au_iu_iu4_t3_t,

   output                    au_iu_iu4_s1_v,
   output [0:`GPR_POOL_ENC-1] au_iu_iu4_s1_a,
   output [0:2]              au_iu_iu4_s1_t,

   output                    au_iu_iu4_s2_v,
   output [0:`GPR_POOL_ENC-1] au_iu_iu4_s2_a,
   output [0:2]              au_iu_iu4_s2_t,

   output                    au_iu_iu4_s3_v,
   output [0:`GPR_POOL_ENC-1] au_iu_iu4_s3_a,
   output [0:2]              au_iu_iu4_s3_t,

   output [0:2]              au_iu_iu4_ilat,
   output                    au_iu_iu4_ord,
   output                    au_iu_iu4_cord,
   output                    au_iu_iu4_spec,
   output                    au_iu_iu4_type_fp,
   output                    au_iu_iu4_type_ap,
   output                    au_iu_iu4_type_spv,
   output                    au_iu_iu4_type_st,
   output                    au_iu_iu4_async_block,

   output                    au_iu_iu4_isload,
   output                    au_iu_iu4_isstore,

   output                    au_iu_iu4_rte_lq,
   output                    au_iu_iu4_rte_sq,
   output                    au_iu_iu4_rte_axu0,
   output                    au_iu_iu4_rte_axu1,

   output                    au_iu_iu4_no_ram,

   //-------------------------------------------------------------------

   output [0:31]             fu_dec_debug
   );

   //------------------------------------------------------------------------------------------------------------------------------------------------------

      wire                      tidn;
      wire                      tiup;

      wire [0:5]                is0_ldst_ra;

      wire [0:7]                iu_au_config_iucr_int;
      wire [0:7]                iu_au_config_iucr_l2;
      wire [0:7]                iu_au_config_iucr_din;
      wire [00:31]              is0_instr;
      wire [0:5]                pri_is0;		// primary opcode
      wire [20:31]              sec_is0;		// secondary opcode
      wire                      av;		// source/target valids
      wire                      bv;
      wire                      cv;
      wire                      tv;
      wire                      isfu_dec_is0;
      wire                      ld_st_is0;
      wire                      isLoad;
      wire                      isStore;

      wire                      st_is0;
      wire                      indexed;
      wire                      fdiv_is0;
      wire                      fsqrt_is0;
      wire                      update_form;
      wire                      forcealign;
      wire                      cr_writer;
      wire                      is0_instr_v;
      wire                      ucode_restart;
      wire                      mffgpr;
      wire                      mftgpr;
      wire                      record_form;
      wire                      fpscr_wr;
      wire                      fpscr_mv;
      wire [0:8]                ldst_tag;
      wire [0:4]                ldst_tag_addr;
      wire                      is0_to_ucode;
      wire                      cordered;
      wire                      ordered;
      wire                      is0_zero_r0;

      wire [0:7]                config_reg_scin;
      wire [0:7]                config_reg_scout;

      wire [0:5]                size;
      wire [3:7]                spare_unused;

      wire                      is0_is_ucode;
      wire                      in_ucode_mode;
      wire                      only_from_ucode;
      wire                      only_graphics_mode;
      wire                      graphics_mode;
      wire                      is0_invalid_kill;
      wire                      is0_invalid_kill_uc;

      wire                      ldst_extpid;
      wire                      single_precision_ldst;
      wire                      int_word_ldst;
      wire                      sign_ext_ldst;
      wire                      io_port;
      wire                      io_port_ext;

      wire                      ignore_flush_is0;

      wire                      is0_kill_or_divsqrt_b;
      wire                      au_iu_is0_i_dec;
      wire                      is0_i_dec_b;
      wire                      no_ram;

      wire                      ram_mode_v;

      wire [0:5]                au_iu_iu4_t1_a6;
      wire [0:5]                au_iu_iu4_t2_a6;
      wire [0:5]                au_iu_iu4_t3_a6;
      wire [0:5]                au_iu_iu4_s1_a6;
      wire [0:5]                au_iu_iu4_s2_a6;
      wire [0:5]                au_iu_iu4_s3_a6;

      // Pervasive
      wire                      pc_iu_func_sl_thold_1;
      wire                      pc_iu_func_sl_thold_0;
      wire                      pc_iu_func_sl_thold_0_b;
      wire                      pc_iu_sg_1;
      wire                      pc_iu_sg_0;
      wire                      force_t;
   //--------------------------------------------------------------

      //-----------------------------------------------
      // pervasive
      //-----------------------------------------------


   tri_plat #(.WIDTH(2)) perv_2to1_reg(
      .vd(vdd),
      .gd(gnd),
      .nclk(nclk),
      .flush(tc_ac_ccflush_dc),
      .din({pc_iu_func_sl_thold_2,pc_iu_sg_2}),
      .q({pc_iu_func_sl_thold_1,pc_iu_sg_1})
   );


   tri_plat #(.WIDTH(2)) perv_1to0_reg(
      .vd(vdd),
      .gd(gnd),
      .nclk(nclk),
      .flush(tc_ac_ccflush_dc),
      .din({pc_iu_func_sl_thold_1,pc_iu_sg_1}),
      .q({pc_iu_func_sl_thold_0,pc_iu_sg_0})
   );


         tri_lcbor  perv_lcbor(
            .clkoff_b(clkoff_b),
            .thold(pc_iu_func_sl_thold_0),
            .sg(pc_iu_sg_0),
            .act_dis(act_dis),
            .force_t(force_t),
            .thold_b(pc_iu_func_sl_thold_0_b)
         );

      assign tidn = 1'b0;
      assign tiup = 1'b1;

      assign is0_instr = iu_au_iu4_instr;
      assign is0_instr_v = iu_au_iu4_instr_v;
      assign ucode_restart = iu_au_ucode_restart;

      assign pri_is0[0:5] = is0_instr[0:5];
      assign sec_is0[20:31] = is0_instr[20:31];

      // update # of inputs and outputs   .i xx   .o xx
      // run "espvhdlexpand iuq_axu_fu_dec.vhdl > iuq_axu_fu_dec_new.vhdl" to regenerate logic below table
      //

      //@@ ESPRESSO TABLE START @@
      // ##################################################################################################
      // .i 18
      // .o 35
      // .ilb pri_is0[0] pri_is0[1] pri_is0[2] pri_is0[3] pri_is0[4] pri_is0[5]
      //      sec_is0[20] sec_is0[21] sec_is0[22] sec_is0[23] sec_is0[24] sec_is0[25] sec_is0[26] sec_is0[27] sec_is0[28] sec_is0[29] sec_is0[30] sec_is0[31]
      // .ob  isfu_dec_is0 tv av bv cv
      //      record_form fpscr_wr cordered ordered fpscr_mv
      //      ld_st_is0 st_is0 indexed update_form forcealign single_precision_ldst int_word_ldst sign_ext_ldst ldst_extpid io_port io_port_ext
      //      size[0] size[1] size[2] size[3] size[4] size[5]
      //      cr_writer mffgpr mftgpr fdiv_is0
      //      fsqrt_is0   only_from_ucode no_ram only_graphics_mode
      // .type fd
      //#
      //#
      // #####################################################################################################################
      //#                                                                       s
      //#                                                                       i
      //#                                                                       n
      //#                                                                       g                                         o
      //#                                                                       l                                         n
      //#                                                                       e                                         l
      //#                                                                       |                                     o   y
      //#                                                                       p                                     n   |
      //#                                                                       r i s                                 l   g
      //#                                                                       e n i                                 y   r
      //#                                                                   u   c t g l  i                            |   a
      //#                                                                   p f i | n d  o                            f   p
      //#                                                                   d o s w | s  |               c            r   h
      //#                                                    f c   f  l     a r i o e t  p     LD/ST     r            o   i
      //#                                                    p o o p  d   i t c o r x | io     size                   m   c
      //#                                                  r s r r s      n e e n d t e or     in        w   mm       | n s
      //#                                                  e c d d c  o s d   a | | | x |t     bytes     r   ff  f    u o |
      //#pri_is0    sec_is0        i                       c r e e r  r t e f l l l l t p|     1to16     i   ft fs    c | m
      //#                          s                       o _ r r _    o x o i d d d p oe     pwrs      t   gg dq    o r o
      //#000000 2 2222222223 3     F      T   A   B   C    r w e e m  s r e r g s s s i rx     oftwo     e   pp ir    d a d
      //#012345 0 1234567890 1     U      V   V   V   V    d r d d v  t e d m n t t t d tt    012345     r   rr vt    e m e
      // #####################################################################################################################

      // 000000 - ---------- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    110011     -   00 00    0 0 0 # reserved
      // 000001 - ---------- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0 # open for vxu new instructions
      // 000010 - ---------- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 000011 - ---------- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 000100 - 000------- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 000100 - 0010------ -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 000100 - 00110000-- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 000100 - 0011000100 -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 000100 - 0011000101 1     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 000100 - 001100011- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 000100 - 0011001--- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 000100 - 001101---- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 000100 - 00111000-- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 000100 - 0011100100 -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 000100 - 0011100101 1     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 000100 - 001110011- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 000100 - 0011101--- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 000100 - 001111---- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 000100 - 01-------- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 000100 - 1--------- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 000101 - ---------- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 000110 - ---------- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 000111 - ---------- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 001--- - ---------- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 010--- - ---------- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 01-0-- - ---------- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 01--0- - ---------- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 01---0 - ---------- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 011111 - 0000000000 -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 011111 1 0000000011 0     0      1   0   0   0    0 0 0 0 -  1 0 1 0 0 0 1 0 0 11    000000     0   10 00    0 0 0 # mfdpx   (DITC to FPR)
      // 011111 1 0000000011 1     0      1   0   0   0    0 0 0 0 -  1 0 1 0 0 0 1 0 0 11    000000     1   10 00    0 0 0 # mfdpx.  (DITC to FPR)
      // 011111 1 0000100011 0     0      1   0   0   0    0 0 0 0 -  1 0 0 0 0 0 1 0 0 10    000000     0   10 00    0 0 0 # mfdp    (DITC to FPR)
      // 011111 1 0000100011 1     0      1   0   0   0    0 0 0 0 -  1 0 0 0 0 0 1 0 0 10    000000     1   10 00    0 0 0 # mfdp.   (DITC to FPR)
      // 011111 1 0001000011 0     0      0   1   0   0    0 0 0 0 -  1 1 1 0 0 0 1 0 0 11    000000     0   01 00    0 0 0 # mtdpx   (DITC from FPR)
      // 011111 1 0001000011 1     0      0   1   0   0    0 0 0 0 -  1 1 1 0 0 0 1 0 0 11    000000     1   01 00    0 0 0 # mtdpx.  (DITC from FPR)
      // 011111 1 0001100011 0     0      0   1   0   0    0 0 0 0 -  1 1 0 0 0 0 1 0 0 10    000000     0   01 00    0 0 0 # mtdp    (DITC from FPR)
      // 011111 1 0001100011 1     0      0   1   0   0    0 0 0 0 -  1 1 0 0 0 0 1 0 0 10    000000     1   01 00    0 0 0 # mtdp.   (DITC from FPR)
      // 011111 - 01-------- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 011111 - 100000---- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 011111 - 10000100-- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 011111 - 100001010- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 011111 - 1000010110 -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 011111 - 1000010111 -     1      1   0   0   0    0 0 0 0 -  1 0 1 0 0 1 0 0 0 00    000100     0   00 00    0 0 0 # lfsx
      // 011111 - 1000011--- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 011111 - 100010---- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 011111 - 10001100-- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 011111 - 100011010- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 011111 - 1000110110 -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 011111 - 1000110111 -     1      1   0   0   0    0 0 0 0 -  1 0 1 1 0 1 0 0 0 00    000100     0   00 00    0 1 0 # lfsux
      // 011111 - 1000111--- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 011111 - 100100---- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 011111 - 10010100-- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 011111 - 100101010- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 011111 - 1001010110 -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 011111 - 1001010111 -     1      1   0   0   0    0 0 0 0 -  1 0 1 0 0 0 0 0 0 00    001000     0   00 00    0 0 0 # lfdx
      // 011111 - 10010110-- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 011111 - 100101110- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 011111 - 1001011110 -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 011111 - 1001011111 -     1      1   0   0   0    0 0 0 0 -  1 0 1 0 0 0 0 0 1 00    001000     0   00 00    0 0 0 # lfdepx
      // 011111 - 100110---- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 011111 - 10011100-- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 011111 - 100111010- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 011111 - 1001110110 -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 011111 - 1001110111 -     1      1   0   0   0    0 0 0 0 -  1 0 1 1 0 0 0 0 0 00    001000     0   00 00    0 1 0 # lfdux
      // 011111 - 1001111100 -     1      1   0   0   0    0 0 0 0 -  1 0 0 0 0 0 1 1 0 00    000000     0   10 00    1 0 1 # mfifgpr (mffgpr for lfiwax)
      // 011111 - 1001111101 -     1      1   0   0   0    0 0 0 0 -  1 0 0 0 0 0 1 0 0 00    000000     0   10 00    1 0 1 # mfixfgpr (mffgpr for lfiwzx)
      // 011111 - 1001111110 -     1      1   0   0   0    0 0 0 0 -  1 0 0 0 0 1 0 0 0 00    000000     0   10 00    1 0 1 # mfsfgpr (mffgpr for lfs, lfsu single)
      // 011111 - 1001111111 -     1      1   0   0   0    0 0 0 0 -  1 0 0 0 0 0 0 0 0 00    000000     0   10 00    1 0 1 # mffgpr (mffgpr for lfd, lfdu double)
      // 011111 - 101000---- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 011111 - 10100100-- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 011111 - 101001010- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 011111 - 1010010110 -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 011111 - 1010010111 -     1      0   1   0   0    0 0 0 0 -  1 1 1 0 0 1 0 0 0 00    000100     0   00 00    0 0 0 # stfsx
      // 011111 - 1010011--- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 011111 - 101010---- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 011111 - 10101100-- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 011111 - 101011010- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 011111 - 1010110110 -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 011111 - 1010110111 -     1      0   1   0   0    0 0 0 0 -  1 1 1 1 0 1 0 0 0 00    000100     0   00 00    0 0 0 # stfsux
      // 011111 - 1010111--- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 011111 - 101100---- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 011111 - 10110100-- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 011111 - 101101010- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 011111 - 1011010110 -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 011111 - 1011010111 -     1      0   1   0   0    0 0 0 0 -  1 1 1 0 0 0 0 0 0 00    001000     0   00 00    0 0 0 # stfdx
      // 011111 - 10110110-- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 011111 - 1011011100 -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 011111 - 1011011101 -     1      0   0   1   0    0 0 0 0 -  1 1 0 0 0 0 1 0 0 00    000000     0   01 00    1 0 1 # mfitgpr (mftgpr for stfiwx integer word)
      // 011111 - 1011011110 -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 011111 - 1011011111 -     1      0   1   0   0    0 0 0 0 -  1 1 1 0 0 0 0 0 1 00    001000     0   00 00    0 0 0 # stfdepx
      // 011111 - 101110---- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 011111 - 10111100-- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 011111 - 101111010- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 011111 - 1011110110 -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 011111 - 1011110111 -     1      0   1   0   0    0 0 0 0 -  1 1 1 1 0 0 0 0 0 00    001000     0   00 00    0 0 0 # stfdux
      // 011111 - 1011111110 -     1      0   0   1   0    0 0 0 0 -  1 1 0 0 0 1 0 0 0 00    000000     0   01 00    1 0 1 # mfstgpr (mftgpr single)
      // 011111 - 1011111111 -     1      0   0   1   0    0 0 0 0 -  1 1 0 0 0 0 0 0 0 00    000000     0   01 00    1 0 1 # mftgpr (mftgpr double)
      // 011111 - 110000---- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 011111 - 11000100-- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 011111 - 110001010- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 011111 - 1100010110 -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      //#011111 - 1100010111 -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0 # lfdpx  (ucoded)
      // 011111 - 1100011--- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 011111 - 11001----- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 011111 - 110100---- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 011111 - 11010100-- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 011111 - 110101010- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 011111 - 1101010110 -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 011111 - 1101010111 -     1      1   0   0   0    0 0 0 0 -  1 0 1 0 0 0 1 1 0 00    000100     0   00 00    0 0 0 # lfiwax
      // 011111 - 1101011--- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 011111 - 1101110111 -     1      1   0   0   0    0 0 0 0 -  1 0 1 0 0 0 1 0 0 00    000100     0   00 00    0 0 0 # lfiwzx
      // 011111 - 111000---- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 011111 - 11100100-- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 011111 - 111001010- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 011111 - 1110010110 -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      //#011111 - 1110010111 -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0 # stfdpx   (ucoded)
      // 011111 - 1110011--- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 011111 - 11101----- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 011111 - 111100---- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 011111 - 11110100-- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 011111 - 111101010- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 011111 - 1111010110 -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 011111 - 1111010111 -     1      0   1   0   0    0 0 0 0 -  1 1 1 0 0 0 1 0 0 00    000100     0   00 00    0 0 0 # stfiwx
      // 011111 - 1111011--- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 011111 - 11111----- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 10---- - ---------- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 110000 - ---------- -     1      1   0   0   0    0 0 0 0 -  1 0 0 0 0 1 0 0 0 00    000100     0   00 00    0 0 0 # lfs
      // 110001 - ---------- -     1      1   0   0   0    0 0 0 0 -  1 0 0 1 0 1 0 0 0 00    000100     0   00 00    0 1 0 # lfsu
      // 110010 - ---------- -     1      1   0   0   0    0 0 0 0 -  1 0 0 0 0 0 0 0 0 00    001000     0   00 00    0 0 0 # lfd
      // 110011 - ---------- -     1      1   0   0   0    0 0 0 0 -  1 0 0 1 0 0 0 0 0 00    001000     0   00 00    0 1 0 # lfdu
      // 110100 - ---------- -     1      0   1   0   0    0 0 0 0 -  1 1 0 0 0 1 0 0 0 00    000100     0   00 00    0 0 0 # stfs
      // 110101 - ---------- -     1      0   1   0   0    0 0 0 0 -  1 1 0 1 0 1 0 0 0 00    000100     0   00 00    0 0 0 # stfsu
      // 110110 - ---------- -     1      0   1   0   0    0 0 0 0 -  1 1 0 0 0 0 0 0 0 00    001000     0   00 00    0 0 0 # stfd
      // 110111 - ---------- -     1      0   1   0   0    0 0 0 0 -  1 1 0 1 0 0 0 0 0 00    001000     0   00 00    0 0 0 # stfdu
      // 111000 - ---------- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      //#111001 - ---------0 0     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0 # lfdp    (ucoded)
      // 111001 - ---------0 1     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111001 - ---------1 -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111010 - ---------- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111011 - 000--0---- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111011 - 0010-0---- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111011 - 00110000-- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111011 - 0011000100 -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111011 - 0011000101 0     1      1   0   1   0    0 0 0 0 -  0 0 0 0 0 - - - 0 00    ------     0   00 00    0 0 1 # fexptes
      // 111011 - 001100011- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111011 - 00110010-- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111011 - 001100110- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111011 - 0011001110 0     0      1   0   1   0    0 0 0 0 -  0 0 0 0 0 0 0 0 0 00    ------     0   00 00    0 0 0 # fcfiwus  (removed)
      // 111011 - 0011001110 1     0      1   0   1   0    1 1 1 0 -  0 0 0 0 0 0 0 0 0 00    ------     1   00 00    0 0 0 # fcfiwus. (removed)
      // 111011 - 0011001111 -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111011 - 00111000-- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111011 - 0011100100 -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111011 - 0011100101 0     1      1   0   1   0    0 0 0 0 -  0 0 0 0 0 - - - 0 00    ------     0   00 00    0 0 1 # floges
      // 111011 - 001110011- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111011 - 0011101--- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111011 - 01---0---- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111011 - 10---0---- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111011 - 1100-0---- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111011 - 1101000--- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111011 - 11010010-- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111011 - 110100110- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111011 - 1101001110 0     1      1   0   1   0    0 1 0 0 -  0 0 0 0 0 0 0 0 0 00    ------     0   00 00    0 0 0 # fcfids
      // 111011 - 1101001110 1     1      1   0   1   0    1 1 1 0 -  0 0 0 0 0 0 0 0 0 00    ------     1   00 00    0 0 0 # fcfids.
      // 111011 - 1101001111 -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111011 - 110110---- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111011 - 1110-0---- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111011 - 1111000--- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111011 - 11110010-- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111011 - 111100110- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111011 - 1111001110 0     1      1   0   1   0    0 1 0 0 -  0 0 0 0 0 0 0 0 0 00    ------     0   00 00    0 0 0 # fcfidus
      // 111011 - 1111001110 1     1      1   0   1   0    1 1 1 0 -  0 0 0 0 0 0 0 0 0 00    ------     1   00 00    0 0 0 # fcfidus.
      // 111011 - 1111001111 -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111011 - 111110---- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111011 - -----10000 -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111011 - -----10001 0     0      1   1   0   1    0 1 1 0 -  0 0 0 0 0 0 0 0 0 00    ------     0   00 00    1 0 0 # fmuls_uc
      // 111011 - -----10001 1     0      1   1   0   1    1 1 1 0 -  0 0 0 0 0 0 0 0 0 00    ------     1   00 00    1 0 0 # fmuls_uc.
      // 111011 - -----10010 0     1      1   1   1   0    0 1 0 1 -  0 0 0 0 0 0 0 0 0 00    ------     0   00 10    0 0 0 # fdivs
      // 111011 - -----10010 1     1      1   1   1   0    1 1 1 1 -  0 0 0 0 0 0 0 0 0 00    ------     1   00 10    0 0 0 # fdivs.
      // 111011 - -----10011 -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111011 - -----10100 0     1      1   1   1   0    0 1 0 0 -  0 0 0 0 0 0 0 0 0 00    ------     0   00 00    0 0 0 # fsubs
      // 111011 - -----10100 1     1      1   1   1   0    1 1 1 0 -  0 0 0 0 0 0 0 0 0 00    ------     1   00 00    0 0 0 # fsubs.
      // 111011 - -----10101 0     1      1   1   1   0    0 1 0 0 -  0 0 0 0 0 0 0 0 0 00    ------     0   00 00    0 0 0 # fadds
      // 111011 - -----10101 1     1      1   1   1   0    1 1 1 0 -  0 0 0 0 0 0 0 0 0 00    ------     1   00 00    0 0 0 # fadds.
      // 111011 - -----10110 0     1      1   0   1   0    0 1 0 1 -  0 0 0 0 0 0 0 0 0 00    ------     0   00 01    0 0 0 # fsqrts
      // 111011 - -----10110 1     1      1   0   1   0    1 1 1 1 -  0 0 0 0 0 0 0 0 0 00    ------     1   00 01    0 0 0 # fsqrts.
      // 111011 - -----10111 -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111011 - -----11000 0     1      1   0   1   0    0 1 0 0 -  0 0 0 0 0 0 0 0 0 00    ------     0   00 00    0 0 0 # fres
      // 111011 - -----11000 1     1      1   0   1   0    1 1 1 0 -  0 0 0 0 0 0 0 0 0 00    ------     1   00 00    0 0 0 # fres.
      // 111011 - -----11001 0     1      1   1   0   1    0 1 0 0 -  0 0 0 0 0 0 0 0 0 00    ------     0   00 00    0 0 0 # fmuls
      // 111011 - -----11001 1     1      1   1   0   1    1 1 1 0 -  0 0 0 0 0 0 0 0 0 00    ------     1   00 00    0 0 0 # fmuls.
      // 111011 - -----11010 0     1      1   0   1   0    0 1 0 0 -  0 0 0 0 0 0 0 0 0 00    ------     0   00 00    0 0 0 # frsqrtes
      // 111011 - -----11010 1     1      1   0   1   0    1 1 1 0 -  0 0 0 0 0 0 0 0 0 00    ------     1   00 00    0 0 0 # frsqrtes.
      // 111011 - -----11011 -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111011 - -----11100 0     1      1   1   1   1    0 1 0 0 -  0 0 0 0 0 0 0 0 0 00    ------     0   00 00    0 0 0 # fmsubs
      // 111011 - -----11100 1     1      1   1   1   1    1 1 1 0 -  0 0 0 0 0 0 0 0 0 00    ------     1   00 00    0 0 0 # fmsubs.
      // 111011 - -----11101 0     1      1   1   1   1    0 1 0 0 -  0 0 0 0 0 0 0 0 0 00    ------     0   00 00    0 0 0 # fmadds
      // 111011 - -----11101 1     1      1   1   1   1    1 1 1 0 -  0 0 0 0 0 0 0 0 0 00    ------     1   00 00    0 0 0 # fmadds.
      // 111011 - -----11110 0     1      1   1   1   1    0 1 0 0 -  0 0 0 0 0 0 0 0 0 00    ------     0   00 00    0 0 0 # fnmsubs
      // 111011 - -----11110 1     1      1   1   1   1    1 1 1 0 -  0 0 0 0 0 0 0 0 0 00    ------     1   00 00    0 0 0 # fnmsubs.
      // 111011 - -----11111 0     1      1   1   1   1    0 1 0 0 -  0 0 0 0 0 0 0 0 0 00    ------     0   00 00    0 0 0 # fnmadds
      // 111011 - -----11111 1     1      1   1   1   1    1 1 1 0 -  0 0 0 0 0 0 0 0 0 00    ------     1   00 00    0 0 0 # fnmadds.
      // 111100 - ---------- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      //#111101 - ---------0 0     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0 # stfdp  (ucoded)
      // 111101 - ---------0 1     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111101 - ---------1 -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111110 - ---------- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      //#111111 - -----1---- -     0                           - - -  0 0             0 00                            0 0 0
      // 111111 - 0000000000 -     1      0   1   1   0    0 1 0 0 -  0 0 0 0 0 0 0 0 0 00    ------     1   00 00    0 0 0 # fcmpu
      // 111111 - 0000000001 -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111111 - 000000001- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111111 - 00000001-- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111111 - 0000001000 0     1      1   1   1   0    0 0 0 0 -  0 0 0 0 0 0 0 0 0 00    ------     0   00 00    0 0 0 # fcpsgn
      // 111111 - 0000001000 1     1      1   1   1   0    1 0 1 0 -  0 0 0 0 0 0 0 0 0 00    ------     1   00 00    0 0 0 # fcpsgn.
      // 111111 - 0000001001 -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111111 - 000000101- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111111 - 0000001100 0     1      1   0   1   0    0 1 0 0 -  0 0 0 0 0 0 0 0 0 00    ------     0   00 00    0 0 0 # frsp
      // 111111 - 0000001100 1     1      1   0   1   0    1 1 1 0 -  0 0 0 0 0 0 0 0 0 00    ------     1   00 00    0 0 0 # frsp.
      // 111111 - 0000001101 -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111111 - 0000001110 0     1      1   0   1   0    0 1 0 0 -  0 0 0 0 0 0 0 0 0 00    ------     0   00 00    0 0 0 # fctiw
      // 111111 - 0000001110 1     1      1   0   1   0    1 1 1 0 -  0 0 0 0 0 0 0 0 0 00    ------     1   00 00    0 0 0 # fctiw.
      // 111111 - 0000001111 0     1      1   0   1   0    0 1 0 0 -  0 0 0 0 0 0 0 0 0 00    ------     0   00 00    0 0 0 # fctiwz
      // 111111 - 0000001111 1     1      1   0   1   0    1 1 1 0 -  0 0 0 0 0 0 0 0 0 00    ------     1   00 00    0 0 0 # fctiwz.
      // 111111 - -----10000 -     1      1   0   1   0    0 0 0 0 -  0 0 0 0 0 0 0 0 0 00    ------     0   00 00    1 0 0 # prenormalization
      // 111111 - -----10001 0     0      1   1   0   1    0 1 1 0 -  0 0 0 0 0 0 0 0 0 00    ------     0   00 00    1 0 0 # fmul_uc
      // 111111 - -----10001 1     0      1   1   0   1    1 1 1 0 -  0 0 0 0 0 0 0 0 0 00    ------     1   00 00    1 0 0 # fmul_uc.
      // 111111 - -----10010 0     1      1   1   1   0    0 1 0 1 -  0 0 0 0 0 0 0 0 0 00    ------     0   00 10    0 0 0 # fdiv
      // 111111 - -----10010 1     1      1   1   1   0    1 1 1 1 -  0 0 0 0 0 0 0 0 0 00    ------     1   00 10    0 0 0 # fdiv.
      // 111111 - -----10011 -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111111 - -----10100 0     1      1   1   1   0    0 1 0 0 -  0 0 0 0 0 0 0 0 0 00    ------     0   00 00    0 0 0 # fsub
      // 111111 - -----10100 1     1      1   1   1   0    1 1 1 0 -  0 0 0 0 0 0 0 0 0 00    ------     1   00 00    0 0 0 # fsub.
      // 111111 - -----10101 0     1      1   1   1   0    0 1 0 0 -  0 0 0 0 0 0 0 0 0 00    ------     0   00 00    0 0 0 # fadd
      // 111111 - -----10101 1     1      1   1   1   0    1 1 1 0 -  0 0 0 0 0 0 0 0 0 00    ------     1   00 00    0 0 0 # fadd.
      // 111111 - -----10110 0     1      1   0   1   0    0 1 0 1 -  0 0 0 0 0 0 0 0 0 00    ------     0   00 01    0 0 0 # fsqrt
      // 111111 - -----10110 1     1      1   0   1   0    1 1 1 1 -  0 0 0 0 0 0 0 0 0 00    ------     1   00 01    0 0 0 # fsqrt.
      // 111111 - -----10111 0     1      1   1   1   1    0 0 0 0 -  0 0 0 0 0 0 0 0 0 00    ------     0   00 00    0 0 0 # fsel
      // 111111 - -----10111 1     1      1   1   1   1    1 0 1 0 -  0 0 0 0 0 0 0 0 0 00    ------     1   00 00    0 0 0 # fsel.
      // 111111 - -----11000 0     1      1   0   1   0    0 1 0 0 -  0 0 0 0 0 0 0 0 0 00    ------     0   00 00    0 0 0 # fre
      // 111111 - -----11000 1     1      1   0   1   0    1 1 1 0 -  0 0 0 0 0 0 0 0 0 00    ------     1   00 00    0 0 0 # fre.
      // 111111 - -----11001 0     1      1   1   0   1    0 1 0 0 -  0 0 0 0 0 0 0 0 0 00    ------     0   00 00    0 0 0 # fmul
      // 111111 - -----11001 1     1      1   1   0   1    1 1 1 0 -  0 0 0 0 0 0 0 0 0 00    ------     1   00 00    0 0 0 # fmul.
      // 111111 - -----11010 0     1      1   0   1   0    0 1 0 0 -  0 0 0 0 0 0 0 0 0 00    ------     0   00 00    0 0 0 # frsqrte
      // 111111 - -----11010 1     1      1   0   1   0    1 1 1 0 -  0 0 0 0 0 0 0 0 0 00    ------     1   00 00    0 0 0 # frsqrte.
      // 111111 - -----11011 -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111111 - -----11100 0     1      1   1   1   1    0 1 0 0 -  0 0 0 0 0 0 0 0 0 00    ------     0   00 00    0 0 0 # fmsub
      // 111111 - -----11100 1     1      1   1   1   1    1 1 1 0 -  0 0 0 0 0 0 0 0 0 00    ------     1   00 00    0 0 0 # fmsub.
      // 111111 - -----11101 0     1      1   1   1   1    0 1 0 0 -  0 0 0 0 0 0 0 0 0 00    ------     0   00 00    0 0 0 # fmadd
      // 111111 - -----11101 1     1      1   1   1   1    1 1 1 0 -  0 0 0 0 0 0 0 0 0 00    ------     1   00 00    0 0 0 # fmadd.
      // 111111 - -----11110 0     1      1   1   1   1    0 1 0 0 -  0 0 0 0 0 0 0 0 0 00    ------     0   00 00    0 0 0 # fnmsub
      // 111111 - -----11110 1     1      1   1   1   1    1 1 1 0 -  0 0 0 0 0 0 0 0 0 00    ------     1   00 00    0 0 0 # fnmsub.
      // 111111 - -----11111 0     1      1   1   1   1    0 1 0 0 -  0 0 0 0 0 0 0 0 0 00    ------     0   00 00    0 0 0 # fnmadd
      // 111111 - -----11111 1     1      1   1   1   1    1 1 1 0 -  0 0 0 0 0 0 0 0 0 00    ------     1   00 00    0 0 0 # fnmadd.
      // 111111 - 0000100000 -     1      0   1   1   0    0 1 0 0 -  0 0 0 0 0 0 0 0 0 00    ------     1   00 00    0 0 0 # fcmpo
      // 111111 - 0000100001 -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111111 - 000010001- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111111 - 000010010- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111111 - 0000100110 0     1      0   0   0   0    0 0 1 0 1  0 0 0 0 0 0 0 0 0 00    ------     0   00 00    0 0 0 # mtfsb1
      // 111111 - 0000100110 1     1      0   0   0   0    1 0 1 0 1  0 0 0 0 0 0 0 0 0 00    ------     1   00 00    0 0 0 # mtfsb1.
      // 111111 - 0000100111 -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111111 - 0000101000 0     1      1   0   1   0    0 0 0 0 -  0 0 0 0 0 0 0 0 0 00    ------     0   00 00    0 0 0 # fneg
      // 111111 - 0000101000 1     1      1   0   1   0    1 0 1 0 -  0 0 0 0 0 0 0 0 0 00    ------     1   00 00    0 0 0 # fneg.
      // 111111 - 0000101001 -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111111 - 000010101- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111111 - 00001011-- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      //#111111 - 000011---- -     0                           - - -  0 0             0 00                            0 0 0
      // 111111 - 0001000000 -     1      0   0   0   0    0 0 1 0 1  0 0 0 0 0 0 0 0 0 00    ------     1   00 00    0 0 0 # mcrfs
      // 111111 - 0001000001 -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111111 - 000100001- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111111 - 000100010- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111111 - 0001000110 0     1      0   0   0   0    0 0 1 0 1  0 0 0 0 0 0 0 0 0 00    ------     0   00 00    0 0 0 # mtfsb0
      // 111111 - 0001000110 1     1      0   0   0   0    1 0 1 0 1  0 0 0 0 0 0 0 0 0 00    ------     1   00 00    0 0 0 # mtfsb0.
      // 111111 - 0001000111 -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111111 - 0001001000 0     1      1   0   1   0    0 0 0 0 -  0 0 0 0 0 0 0 0 0 00    ------     0   00 00    0 0 0 # fmr
      // 111111 - 0001001000 1     1      1   0   1   0    1 0 1 0 -  0 0 0 0 0 0 0 0 0 00    ------     1   00 00    0 0 0 # fmr.
      // 111111 - 0001001001 -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111111 - 000100101- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111111 - 00010011-- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      //#111111 - 000101---- -     0                           - - -  0 0             0 00                            0 0 0
      // 111111 - 000110---- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      //#111111 - 000111---- -     0                           - - -  0 0             0 00                            0 0 0
      // 111111 - 0010000000 -     1      0   1   1   0    0 0 0 0 -  0 0 0 0 0 0 0 0 0 00    ------     1   00 00    0 0 0 # ftdiv
      // 111111 - 001000010- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111111 - 0010000110 0     1      0   0   0   0    0 0 1 0 1  0 0 0 0 0 0 0 0 0 00    ------     0   00 00    0 0 0 # mtfsfi
      // 111111 - 0010000110 1     1      0   0   0   0    1 0 1 0 1  0 0 0 0 0 0 0 0 0 00    ------     1   00 00    0 0 0 # mtfsfi.
      // 111111 - 0010000111 -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111111 - 0010001000 0     1      1   0   1   0    0 0 0 0 -  0 0 0 0 0 0 0 0 0 00    ------     0   00 00    0 0 0 # fnabs
      // 111111 - 0010001000 1     1      1   0   1   0    1 0 1 0 -  0 0 0 0 0 0 0 0 0 00    ------     1   00 00    0 0 0 # fnabs.
      // 111111 - 0010001001 -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111111 - 001000101- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111111 - 001000110- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111111 - 0010001110 0     1      1   0   1   0    0 1 0 0 -  0 0 0 0 0 0 0 0 0 00    ------     0   00 00    0 0 0 # fctiwu
      // 111111 - 0010001110 1     1      1   0   1   0    1 1 1 0 -  0 0 0 0 0 0 0 0 0 00    ------     1   00 00    0 0 0 # fctiwu.
      // 111111 - 0010001111 0     1      1   0   1   0    0 1 0 0 -  0 0 0 0 0 0 0 0 0 00    ------     0   00 00    0 0 0 # fctiduz
      // 111111 - 0010001111 1     1      1   0   1   0    1 1 1 0 -  0 0 0 0 0 0 0 0 0 00    ------     1   00 00    0 0 0 # fctiduz.
      //#111111 - 001001---- -     0                           - - -  0 0             0 00                            0 0 0
      // 111111 - 0010100000 -     1      0   0   1   0    0 0 0 0 -  0 0 0 0 0 0 0 0 0 00    ------     1   00 00    0 0 0 # ftsqrt
      //#111111 - 001011---- -     0                           - - -  0 0             0 00                            0 0 0
      // 111111 - 0011000--- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111111 - 00110010-- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111111 - 001100110- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111111 - 0011001110 0     0      1   0   1   0    0 1 0 0 -  0 0 0 0 0 0 0 0 0 00    ------     0   00 00    0 0 0 # fcfiwu  (removed)
      // 111111 - 0011001110 1     0      1   0   1   0    1 1 1 0 -  0 0 0 0 0 0 0 0 0 00    ------     1   00 00    0 0 0 # fcfiwu. (removed)
      // 111111 - 0011001111 -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      //#111111 - 001101---- -     0                           - - -  0 0             0 00                            0 0 0
      // 111111 - 001110---- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      //#111111 - 001111---- -     0                           - - -  0 0             0 00                            0 0 0
      // 111111 - 0100000--- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111111 - 0100001000 0     1      1   0   1   0    0 0 0 0 -  0 0 0 0 0 0 0 0 0 00    ------     0   00 00    0 0 0 # fabs
      // 111111 - 0100001000 1     1      1   0   1   0    1 0 1 0 -  0 0 0 0 0 0 0 0 0 00    ------     1   00 00    0 0 0 # fabs.
      // 111111 - 0100001001 -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111111 - 010000101- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111111 - 01000011-- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      //#111111 - 010001---- -     0                           - - -  0 0             0 00                            0 0 0
      // 111111 - 010010---- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      //#111111 - 010011---- -     0                           - - -  0 0             0 00                            0 0 0
      // 111111 - 010100---- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      //#111111 - 010101---- -     0                           - - -  0 0             0 00                            0 0 0
      // 111111 - 010110---- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      //#111111 - 010111---- -     0                           - - -  0 0             0 00                            0 0 0
      // 111111 - 0110000--- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111111 - 0110001000 0     1      1   0   1   0    0 1 0 0 -  0 0 0 0 0 0 0 0 0 00    ------     0   00 00    0 0 0 # frin
      // 111111 - 0110001000 1     1      1   0   1   0    1 1 1 0 -  0 0 0 0 0 0 0 0 0 00    ------     1   00 00    0 0 0 # frin.
      // 111111 - 0110001001 -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111111 - 011000101- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111111 - 01100011-- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      //#111111 - 011001---- -     0                           - - -  0 0   0         0 00                            0 0 0
      // 111111 - 0110100--- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111111 - 0110101000 0     1      1   0   1   0    0 1 0 0 -  0 0 0 0 0 0 0 0 0 00    ------     0   00 00    0 0 0 # friz
      // 111111 - 0110101000 1     1      1   0   1   0    1 1 1 0 -  0 0 0 0 0 0 0 0 0 00    ------     1   00 00    0 0 0 # friz.
      // 111111 - 0110101001 -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111111 - 011010101- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111111 - 01101011-- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      //#111111 - 011011---- -     0                           - - -  0 0   0         0 00                            0 0 0
      // 111111 - 0111000--- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111111 - 0111001000 0     1      1   0   1   0    0 1 0 0 -  0 0 0 0 0 0 0 0 0 00    ------     0   00 00    0 0 0 # frip
      // 111111 - 0111001000 1     1      1   0   1   0    1 1 1 0 -  0 0 0 0 0 0 0 0 0 00    ------     1   00 00    0 0 0 # frip.
      // 111111 - 0111001001 -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111111 - 011100101- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111111 - 01110011-- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      //#111111 - 011101---- -     0                           - - -  0 0   0         0 00                            0 0 0
      // 111111 - 0111100--- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111111 - 0111101000 0     1      1   0   1   0    0 1 0 0 -  0 0 0 0 0 0 0 0 0 00    ------     0   00 00    0 0 0 # frim
      // 111111 - 0111101000 1     1      1   0   1   0    1 1 1 0 -  0 0 0 0 0 0 0 0 0 00    ------     1   00 00    0 0 0 # frim.
      // 111111 - 0111101001 -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111111 - 011110101- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111111 - 01111011-- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      //#111111 - 011111---- -     0                           - - -  0 0             0 00                            0 0 0
      // 111111 - 100000---- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      //#111111 - 100001---- -     0                           - - -  0 0             0 00                            0 0 0
      // 111111 - 100010---- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      //#111111 - 100011---- -     0                           - - -  0 0             0 00                            0 0 0
      // 111111 - 10010000-- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111111 - 100100010- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111111 - 1001000110 -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111111 - 1001000111 0     1      1   0   0   0    0 0 1 0 -  0 0 0 0 0 0 0 0 0 00    ------     0   00 00    0 0 0 # mffs
      // 111111 - 1001000111 1     1      1   0   0   0    1 0 1 0 -  0 0 0 0 0 0 0 0 0 00    ------     1   00 00    0 0 0 # mffs.
      // 111111 - 1001001--- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      //#111111 - 100101---- -     0                           - - -  0 0             0 00                            0 0 0
      // 111111 - 100110---- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      //#111111 - 100111---- -     0                           - - -  0 0             0 00                            0 0 0
      // 111111 - 101000---- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      //#111111 - 101001---- -     0                           - - -  0 0             0 00                            0 0 0
      // 111111 - 101010---- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      //#111111 - 101011---- -     0                           - - -  0 0             0 00                            0 0 0
      // 111111 - 10110000-- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111111 - 101100010- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111111 - 1011000110 -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111111 - 1011000111 0     1      0   0   1   0    0 0 1 0 1  0 0 0 0 0 0 0 0 0 00    ------     0   00 00    0 0 0 # mtfsf
      // 111111 - 1011000111 1     1      0   0   1   0    1 0 1 0 1  0 0 0 0 0 0 0 0 0 00    ------     1   00 00    0 0 0 # mtfsf.
      // 111111 - 1011001--- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      //#111111 - 101101---- -     0                           - - -  0 0             0 00                            0 0 0
      // 111111 - 101110---- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      //#111111 - 101111---- -     0                           - - -  0 0             0 00                            0 0 0
      // 111111 - 110000---- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      //#111111 - 110001---- -     0                           - - -  0 0             0 00                            0 0 0
      // 111111 - 1100100--- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111111 - 11001010-- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111111 - 110010110- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111111 - 1100101110 0     1      1   0   1   0    0 1 0 0 -  0 0 0 0 0 0 0 0 0 00    ------     0   00 00    0 0 0 # fctid
      // 111111 - 1100101110 1     1      1   0   1   0    1 1 1 0 -  0 0 0 0 0 0 0 0 0 00    ------     1   00 00    0 0 0 # fctid.
      // 111111 - 1100101111 0     1      1   0   1   0    0 1 0 0 -  0 0 0 0 0 0 0 0 0 00    ------     0   00 00    0 0 0 # fctidz
      // 111111 - 1100101111 1     1      1   0   1   0    1 1 1 0 -  0 0 0 0 0 0 0 0 0 00    ------     1   00 00    0 0 0 # fctidz.

      //#111111 - 110011---- -     0                           - - -  0 0             0 00                            0 0 0
      // 111111 - 1101000--- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111111 - 11010010-- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111111 - 110100110- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111111 - 1101001110 0     1      1   0   1   0    0 1 0 0 -  0 0 0 0 0 0 0 0 0 00    ------     0   00 00    0 0 0 # fcfid
      // 111111 - 1101001110 1     1      1   0   1   0    1 1 1 0 -  0 0 0 0 0 0 0 0 0 00    ------     1   00 00    0 0 0 # fcfid.
      // 111111 - 1101001111 -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      //#111111 - 110101---- -     0                           - - -  0 0             0 00                            0 0 0
      // 111111 - 110110---- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      //#111111 - 110111---- -     0                           - - -  0 0             0 00                            0 0 0
      // 111111 - 111000---- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      //#111111 - 111001---- -     0                           - - -  0 0             0 00                            0 0 0
      // 111111 - 1110100--- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111111 - 11101010-- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111111 - 111010110- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    ------     -   00 00    0 0 0
      // 111111 - 1110101110 0     1      1   0   1   0    0 1 0 0 -  0 0 0 0 0 0 0 0 0 00    ------     0   00 00    0 0 0 # fctidu
      // 111111 - 1110101110 1     1      1   0   1   0    1 1 1 0 -  0 0 0 0 0 0 0 0 0 00    ------     1   00 00    0 0 0 # fctidu.
      // 111111 - 1110101111 0     1      1   0   1   0    0 1 0 0 -  0 0 0 0 0 0 0 0 0 00    ------     0   00 00    0 0 0 # fctiwuz
      // 111111 - 1110101111 1     1      1   0   1   0    1 1 1 0 -  0 0 0 0 0 0 0 0 0 00    ------     1   00 00    0 0 0 # fctiwuz.
      //#111111 - 111011---- -     0                           - - -  0 0             0 00                            0 0 0
      // 111111 - 1111000--- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    000000     -   00 00    0 0 0
      // 111111 - 11110010-- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    000000     -   00 00    0 0 0
      // 111111 - 111100110- -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    000000     -   00 00    0 0 0
      // 111111 - 1111001110 0     1      1   0   1   0    0 1 0 0 -  0 0 0 0 0 0 0 0 0 00    ------     0   00 00    0 0 0 # fcfidu
      // 111111 - 1111001110 1     1      1   0   1   0    1 1 1 0 -  0 0 0 0 0 0 0 0 0 00    ------     1   00 00    0 0 0 # fcfidu.
      // 111111 - 1111001111 -     0      -   -   -   -    - - - - -  0 0 - 0 - - - - 0 00    000000     -   00 00    0 0 0
      //#111111 - 111101---- -     0                           - - -  0 0             0 00                            0 0 0
      //#111111 - 111110---- -     0      -   -   -   -    - - - - -  0 0 - 0 1 0 0 0 0 00    ------     -   00 00    1 0 0 # reserve for
      // 111111 - 111111---- -     0      -   -   -   -    - - - - -  - - - - 1 - - - - --    110011     -   -- --    - - - # no more <=0

      // #########################################################################
      // .e
      //@@ ESPRESSO TABLE END @@

//@@ ESPRESSO LOGIC START @@
// logic generated on: Tue May  3 12:09:00 2011
assign isfu_dec_is0 =  ( pri_is0[0] &  pri_is0[1] &  pri_is0[3] &  pri_is0[4]
		 &  pri_is0[5] & ~sec_is0[21] & ~sec_is0[22]
		 & ~sec_is0[23] & ~sec_is0[24] & ~sec_is0[25]
		 &  sec_is0[27] & ~sec_is0[29] & ~sec_is0[30]) |
		( pri_is0[0] &  pri_is0[1] & ~pri_is0[3] &  pri_is0[4]
		 &  pri_is0[5] & ~sec_is0[21] & ~sec_is0[22]
		 &  sec_is0[23] &  sec_is0[24] & ~sec_is0[27]
		 &  sec_is0[28] & ~sec_is0[29] &  sec_is0[30]
		 & ~sec_is0[31]) |
		( pri_is0[0] &  pri_is0[1] &  pri_is0[3] &  pri_is0[4]
		 &  pri_is0[5] & ~sec_is0[21] &  sec_is0[22]
		 &  sec_is0[23] &  sec_is0[27] & ~sec_is0[28]
		 & ~sec_is0[29] & ~sec_is0[30]) |
		( pri_is0[1] &  pri_is0[2] &  pri_is0[3] &  pri_is0[4]
		 &  pri_is0[5] &  sec_is0[21] & ~sec_is0[23]
		 &  sec_is0[24] &  sec_is0[26] & ~sec_is0[27]
		 &  sec_is0[28] &  sec_is0[29] &  sec_is0[30]) |
		( pri_is0[0] &  pri_is0[1] &  pri_is0[4] &  pri_is0[5]
		 &  sec_is0[21] &  sec_is0[22] &  sec_is0[24]
		 & ~sec_is0[25] &  sec_is0[27] &  sec_is0[28]
		 &  sec_is0[29] & ~sec_is0[30]) |
		( pri_is0[1] &  pri_is0[2] &  pri_is0[3] &  pri_is0[4]
		 &  pri_is0[5] &  sec_is0[21] &  sec_is0[24]
		 & ~sec_is0[25] &  sec_is0[26] & ~sec_is0[27]
		 &  sec_is0[28] &  sec_is0[29] &  sec_is0[30]) |
		( pri_is0[1] &  pri_is0[2] &  pri_is0[3] &  pri_is0[4]
		 &  pri_is0[5] &  sec_is0[21] & ~sec_is0[22]
		 &  sec_is0[26] & ~sec_is0[27] &  sec_is0[28]
		 &  sec_is0[29] &  sec_is0[30]) |
		( pri_is0[0] &  pri_is0[1] &  pri_is0[3] &  pri_is0[4]
		 &  pri_is0[5] & ~sec_is0[21] & ~sec_is0[24]
		 & ~sec_is0[25] &  sec_is0[27] & ~sec_is0[28]
		 & ~sec_is0[29] & ~sec_is0[30]) |
		( pri_is0[0] &  pri_is0[1] &  pri_is0[3] &  pri_is0[4]
		 &  pri_is0[5] & ~sec_is0[21] & ~sec_is0[22]
		 & ~sec_is0[23] & ~sec_is0[24] & ~sec_is0[28]
		 & ~sec_is0[29] & ~sec_is0[30]) |
		( pri_is0[0] &  pri_is0[1] &  pri_is0[3] &  pri_is0[4]
		 &  pri_is0[5] &  sec_is0[21] &  sec_is0[22]
		 & ~sec_is0[24] &  sec_is0[25] &  sec_is0[27]
		 &  sec_is0[28] &  sec_is0[29]) |
		( pri_is0[1] &  pri_is0[2] &  pri_is0[3] &  pri_is0[4]
		 &  pri_is0[5] &  sec_is0[21] & ~sec_is0[22]
		 & ~sec_is0[23] &  sec_is0[24] &  sec_is0[25]
		 &  sec_is0[26] &  sec_is0[27] &  sec_is0[28]) |
		( pri_is0[0] &  pri_is0[1] &  pri_is0[3] &  pri_is0[4]
		 &  pri_is0[5] &  sec_is0[21] & ~sec_is0[22]
		 &  sec_is0[24] & ~sec_is0[25] & ~sec_is0[27]
		 &  sec_is0[28] &  sec_is0[29] &  sec_is0[30]) |
		( pri_is0[0] &  pri_is0[1] &  pri_is0[3] &  pri_is0[4]
		 &  pri_is0[5] & ~sec_is0[21] & ~sec_is0[22]
		 & ~sec_is0[23] & ~sec_is0[25] & ~sec_is0[28]
		 & ~sec_is0[29] & ~sec_is0[30]) |
		( pri_is0[1] &  pri_is0[2] &  pri_is0[3] &  pri_is0[4]
		 &  pri_is0[5] &  sec_is0[21] & ~sec_is0[22]
		 &  sec_is0[24] &  sec_is0[26] &  sec_is0[28]
		 &  sec_is0[29] &  sec_is0[30]) |
		( pri_is0[1] &  pri_is0[2] &  pri_is0[3] &  pri_is0[4]
		 &  pri_is0[5] &  sec_is0[21] & ~sec_is0[22]
		 &  sec_is0[23] &  sec_is0[24] & ~sec_is0[25]
		 &  sec_is0[26] &  sec_is0[27] &  sec_is0[28]
		 &  sec_is0[30]) |
		( pri_is0[0] &  pri_is0[1] &  pri_is0[3] &  pri_is0[4]
		 &  pri_is0[5] & ~sec_is0[21] & ~sec_is0[22]
		 & ~sec_is0[23] & ~sec_is0[24] &  sec_is0[25]
		 & ~sec_is0[27] &  sec_is0[28] &  sec_is0[29]
		 & ~sec_is0[30]) |
		( pri_is0[0] &  pri_is0[1] &  pri_is0[3] &  pri_is0[4]
		 &  pri_is0[5] & ~sec_is0[21] & ~sec_is0[22]
		 & ~sec_is0[24] & ~sec_is0[27] & ~sec_is0[28]
		 & ~sec_is0[29] & ~sec_is0[30]) |
		( pri_is0[0] &  pri_is0[1] &  pri_is0[3] &  pri_is0[4]
		 &  pri_is0[5] & ~sec_is0[21] & ~sec_is0[22]
		 &  sec_is0[23] & ~sec_is0[24] & ~sec_is0[25]
		 &  sec_is0[28] &  sec_is0[29] & ~sec_is0[30]) |
		( pri_is0[0] &  pri_is0[1] &  pri_is0[3] &  pri_is0[4]
		 &  pri_is0[5] & ~sec_is0[21] & ~sec_is0[22]
		 & ~sec_is0[23] &  sec_is0[24] & ~sec_is0[25]
		 & ~sec_is0[27] &  sec_is0[28] &  sec_is0[29]
		 & ~sec_is0[30]) |
		( pri_is0[0] &  pri_is0[1] &  pri_is0[3] &  pri_is0[4]
		 &  pri_is0[5] & ~sec_is0[21] & ~sec_is0[22]
		 & ~sec_is0[24] & ~sec_is0[25] &  sec_is0[27]
		 &  sec_is0[28] &  sec_is0[29]) |
		( pri_is0[1] &  pri_is0[2] &  pri_is0[3] &  pri_is0[4]
		 &  pri_is0[5] &  sec_is0[21] & ~sec_is0[22]
		 &  sec_is0[24] &  sec_is0[25] &  sec_is0[26]
		 &  sec_is0[27] &  sec_is0[28] &  sec_is0[29]) |
		( pri_is0[0] &  pri_is0[1] &  pri_is0[4] &  pri_is0[5]
		 &  sec_is0[26] &  sec_is0[27] & ~sec_is0[29]) |
		( pri_is0[0] &  pri_is0[1] &  pri_is0[4] &  pri_is0[5]
		 &  sec_is0[26] &  sec_is0[29] & ~sec_is0[30]) |
		( pri_is0[0] &  pri_is0[1] &  pri_is0[4] &  pri_is0[5]
		 &  sec_is0[26] &  sec_is0[28] & ~sec_is0[29]) |
		( pri_is0[0] &  pri_is0[1] &  pri_is0[4] &  pri_is0[5]
		 &  sec_is0[26] &  sec_is0[27] &  sec_is0[28]) |
		( pri_is0[0] &  pri_is0[1] & ~pri_is0[2]) |
		( pri_is0[0] &  pri_is0[1] &  pri_is0[3] &  pri_is0[4]
		 &  pri_is0[5] &  sec_is0[26] &  sec_is0[28]) |
		( pri_is0[0] &  pri_is0[1] &  pri_is0[3] &  pri_is0[4]
		 &  pri_is0[5] &  sec_is0[26] & ~sec_is0[30]);

assign tv =  (~pri_is0[3] &  sec_is0[30] & ~sec_is0[31]) |
	( pri_is0[2] &  pri_is0[4] & ~sec_is0[21] &  sec_is0[22]) |
	( pri_is0[2] &  sec_is0[20] & ~sec_is0[23] & ~sec_is0[24]
	 & ~sec_is0[26] & ~sec_is0[27] & ~sec_is0[28] &  sec_is0[29]
	 &  sec_is0[30]) |
	( pri_is0[2] &  sec_is0[22] & ~sec_is0[23] &  sec_is0[24]
	 &  sec_is0[26] & ~sec_is0[27] &  sec_is0[28] &  sec_is0[29]
	 &  sec_is0[30]) |
	( pri_is0[2] &  pri_is0[4] &  sec_is0[22] & ~sec_is0[24]
	 &  sec_is0[27]) |
	( pri_is0[2] &  pri_is0[4] &  sec_is0[21] & ~sec_is0[22]
	 & ~sec_is0[23] &  sec_is0[28]) |
	( pri_is0[0] &  pri_is0[2] &  pri_is0[4] & ~sec_is0[25]
	 &  sec_is0[27]) |
	( pri_is0[0] &  pri_is0[2] &  pri_is0[4] & ~sec_is0[23]
	 &  sec_is0[27]) |
	( pri_is0[0] &  pri_is0[2] &  pri_is0[4] &  sec_is0[26]) |
	(~pri_is0[2] & ~pri_is0[3]);

assign av =  ( pri_is0[3] &  sec_is0[20] & ~sec_is0[22] & ~sec_is0[23]
	 &  sec_is0[24] & ~sec_is0[26] & ~sec_is0[27] & ~sec_is0[28]
	 &  sec_is0[29] &  sec_is0[30]) |
	( pri_is0[0] &  pri_is0[3] &  pri_is0[4] & ~sec_is0[22]
	 & ~sec_is0[23] & ~sec_is0[24] & ~sec_is0[25] & ~sec_is0[26]
	 & ~sec_is0[28]) |
	( pri_is0[0] &  pri_is0[3] &  pri_is0[4] & ~sec_is0[23]
	 &  sec_is0[25] & ~sec_is0[26] & ~sec_is0[27] & ~sec_is0[29]) |
	(~pri_is0[0] &  sec_is0[21] &  sec_is0[23] &  sec_is0[24]
	 & ~sec_is0[25] &  sec_is0[29]) |
	( pri_is0[0] &  pri_is0[3] &  pri_is0[4] & ~sec_is0[24]
	 & ~sec_is0[25] & ~sec_is0[26] & ~sec_is0[27] & ~sec_is0[29]
	 & ~sec_is0[30]) |
	(~pri_is0[0] &  sec_is0[21] & ~sec_is0[22] &  sec_is0[23]
	 & ~sec_is0[27]) |
	( pri_is0[0] &  pri_is0[2] &  pri_is0[4] &  sec_is0[26]
	 &  sec_is0[27] &  sec_is0[28]) |
	( pri_is0[0] &  pri_is0[2] &  pri_is0[4] &  sec_is0[26]
	 & ~sec_is0[27] & ~sec_is0[28] &  sec_is0[29]) |
	( pri_is0[0] &  pri_is0[2] &  pri_is0[4] &  sec_is0[26]
	 &  sec_is0[28] & ~sec_is0[29]) |
	( pri_is0[0] &  pri_is0[2] &  sec_is0[26] &  sec_is0[30]) |
	( pri_is0[1] & ~pri_is0[2] &  pri_is0[3]);

assign bv =  (~pri_is0[0] &  sec_is0[21] & ~sec_is0[25] & ~sec_is0[29]) |
	( pri_is0[2] & ~pri_is0[3] &  sec_is0[28] &  sec_is0[30]
	 & ~sec_is0[31]) |
	(~pri_is0[0] &  sec_is0[21] &  sec_is0[23] &  sec_is0[25]
	 &  sec_is0[27] &  sec_is0[28] &  sec_is0[29]) |
	( pri_is0[0] &  pri_is0[2] &  pri_is0[4] & ~sec_is0[24]
	 & ~sec_is0[27] & ~sec_is0[28] & ~sec_is0[29] & ~sec_is0[30]) |
	( pri_is0[2] &  pri_is0[4] &  sec_is0[22] & ~sec_is0[24]
	 & ~sec_is0[26]) |
	( pri_is0[0] &  pri_is0[2] &  pri_is0[4] &  sec_is0[23]
	 &  sec_is0[24] & ~sec_is0[25] &  sec_is0[29]) |
	( pri_is0[0] &  pri_is0[2] &  pri_is0[4] & ~sec_is0[25]
	 & ~sec_is0[26] &  sec_is0[27]) |
	( pri_is0[0] &  pri_is0[2] &  pri_is0[4] & ~sec_is0[21]
	 &  sec_is0[24] &  sec_is0[27] & ~sec_is0[30]) |
	( pri_is0[0] &  pri_is0[2] &  sec_is0[26] &  sec_is0[28]
	 &  sec_is0[30]) |
	( pri_is0[0] &  pri_is0[2] &  pri_is0[4] & ~sec_is0[23]
	 & ~sec_is0[26] &  sec_is0[27]) |
	( pri_is0[0] &  pri_is0[2] &  pri_is0[4] &  sec_is0[26]
	 & ~sec_is0[30]);

assign cv =  ( pri_is0[0] &  pri_is0[2] &  sec_is0[26] & ~sec_is0[28]
	 &  sec_is0[30]) |
	( pri_is0[0] &  pri_is0[2] &  sec_is0[26] &  sec_is0[29]
	 &  sec_is0[30]) |
	( pri_is0[0] &  pri_is0[2] &  pri_is0[4] &  sec_is0[26]
	 &  sec_is0[27] &  sec_is0[28]);

assign record_form =  ( pri_is0[0] &  pri_is0[2] & ~sec_is0[21] &  sec_is0[24]
	 &  sec_is0[27] &  sec_is0[31]) |
		( pri_is0[0] &  pri_is0[2] & ~sec_is0[23] &  sec_is0[29]
		 &  sec_is0[31]) |
		( pri_is0[0] &  pri_is0[2] & ~sec_is0[25] &  sec_is0[28]
		 &  sec_is0[29] &  sec_is0[31]) |
		( pri_is0[2] &  sec_is0[22] & ~sec_is0[24]
		 &  sec_is0[27] &  sec_is0[31]) |
		( pri_is0[0] &  pri_is0[2] & ~sec_is0[23] &  sec_is0[27]
		 &  sec_is0[31]) |
		( pri_is0[0] &  pri_is0[2] & ~sec_is0[25] &  sec_is0[27]
		 &  sec_is0[31]) |
		( pri_is0[0] &  pri_is0[2] &  sec_is0[26] &  sec_is0[30]
		 &  sec_is0[31]) |
		( pri_is0[0] &  pri_is0[2] &  sec_is0[26] &  sec_is0[29]
		 &  sec_is0[31]) |
		( pri_is0[0] &  pri_is0[2] &  sec_is0[26] &  sec_is0[28]
		 &  sec_is0[31]) |
		( pri_is0[0] &  pri_is0[2] &  sec_is0[26] &  sec_is0[27]
		 &  sec_is0[31]);

assign fpscr_wr =  ( pri_is0[2] & ~pri_is0[3] & ~sec_is0[30] &  sec_is0[31]) |
	( pri_is0[0] &  pri_is0[2] &  pri_is0[4] & ~sec_is0[23]
	 & ~sec_is0[24] & ~sec_is0[26] & ~sec_is0[27] & ~sec_is0[29]) |
	( pri_is0[2] &  pri_is0[4] &  sec_is0[22] & ~sec_is0[25]
	 &  sec_is0[27] &  sec_is0[29]) |
	( pri_is0[2] &  pri_is0[4] &  sec_is0[21] & ~sec_is0[24]
	 &  sec_is0[27]) |
	( pri_is0[2] &  pri_is0[4] & ~sec_is0[21] &  sec_is0[22]
	 &  sec_is0[23] &  sec_is0[27]) |
	( pri_is0[0] &  pri_is0[2] &  sec_is0[26] & ~sec_is0[29]
	 &  sec_is0[30]) |
	( pri_is0[0] &  pri_is0[2] &  pri_is0[4] &  sec_is0[26]
	 &  sec_is0[28] & ~sec_is0[30]) |
	( pri_is0[0] &  pri_is0[2] &  pri_is0[3] &  pri_is0[4]
	 & ~sec_is0[25] &  sec_is0[27] &  sec_is0[28]) |
	( pri_is0[0] &  pri_is0[2] &  pri_is0[4] &  sec_is0[26]
	 &  sec_is0[29] & ~sec_is0[30]) |
	( pri_is0[0] &  pri_is0[2] &  pri_is0[4] &  sec_is0[26]
	 &  sec_is0[27]);

assign cordered =  ( pri_is0[2] & ~sec_is0[21] &  sec_is0[22] &  sec_is0[27]
	 &  sec_is0[31]) |
	( pri_is0[0] &  pri_is0[2] &  pri_is0[4] & ~sec_is0[23]
	 &  sec_is0[24] & ~sec_is0[26] & ~sec_is0[27]) |
	( pri_is0[0] &  pri_is0[2] &  pri_is0[4] & ~sec_is0[23]
	 & ~sec_is0[26] & ~sec_is0[27] &  sec_is0[29]) |
	( pri_is0[2] &  sec_is0[22] & ~sec_is0[24] &  sec_is0[27]
	 &  sec_is0[31]) |
	( pri_is0[0] &  pri_is0[2] &  pri_is0[4] & ~sec_is0[25]
	 & ~sec_is0[26] & ~sec_is0[27] &  sec_is0[28] &  sec_is0[29]) |
	( pri_is0[0] &  pri_is0[2] & ~sec_is0[23] &  sec_is0[27]
	 &  sec_is0[31]) |
	( pri_is0[0] &  pri_is0[2] & ~sec_is0[25] &  sec_is0[27]
	 &  sec_is0[31]) |
	( pri_is0[0] &  pri_is0[2] &  sec_is0[26] & ~sec_is0[27]
	 & ~sec_is0[28] &  sec_is0[30]) |
	( pri_is0[0] &  pri_is0[2] &  sec_is0[26] &  sec_is0[29]
	 &  sec_is0[31]) |
	( pri_is0[0] &  pri_is0[2] &  sec_is0[26] &  sec_is0[27]
	 &  sec_is0[31]) |
	( pri_is0[0] &  pri_is0[2] &  sec_is0[26] &  sec_is0[28]
	 &  sec_is0[31]);

assign ordered =  ( pri_is0[0] &  pri_is0[2] &  pri_is0[4] &  sec_is0[26]
	 & ~sec_is0[27] &  sec_is0[29] & ~sec_is0[30]);

assign fpscr_mv =  ( pri_is0[0] &  pri_is0[4] & ~sec_is0[25] &  sec_is0[28]
	 &  sec_is0[29]) |
	( pri_is0[0] &  pri_is0[4] & ~sec_is0[23]);

assign ld_st_is0 =  (~pri_is0[0] &  pri_is0[1] &  pri_is0[2] &  pri_is0[3]
	 &  pri_is0[4] &  pri_is0[5] &  sec_is0[20] & ~sec_is0[21]
	 & ~sec_is0[22] & ~sec_is0[23] & ~sec_is0[26] & ~sec_is0[27]
	 & ~sec_is0[28] &  sec_is0[29] &  sec_is0[30]) |
		(~pri_is0[0] &  pri_is0[1] &  pri_is0[2] &  pri_is0[3]
		 &  pri_is0[4] &  pri_is0[5] &  sec_is0[21]
		 & ~sec_is0[22] & ~sec_is0[23] &  sec_is0[24]
		 &  sec_is0[25] &  sec_is0[26] &  sec_is0[27]
		 &  sec_is0[28]) |
		(~pri_is0[0] &  pri_is0[1] &  pri_is0[2] &  pri_is0[3]
		 &  pri_is0[4] &  pri_is0[5] &  sec_is0[21]
		 & ~sec_is0[22] &  sec_is0[23] &  sec_is0[24]
		 & ~sec_is0[25] &  sec_is0[26] &  sec_is0[27]
		 &  sec_is0[28] &  sec_is0[30]) |
		(~pri_is0[0] &  pri_is0[1] &  pri_is0[2] &  pri_is0[3]
		 &  pri_is0[4] &  pri_is0[5] &  sec_is0[21]
		 & ~sec_is0[22] &  sec_is0[24] &  sec_is0[25]
		 &  sec_is0[26] &  sec_is0[27] &  sec_is0[28]
		 &  sec_is0[29]) |
		(~pri_is0[0] &  pri_is0[1] &  pri_is0[2] &  pri_is0[3]
		 &  pri_is0[4] &  pri_is0[5] &  sec_is0[21]
		 &  sec_is0[24] & ~sec_is0[25] &  sec_is0[26]
		 & ~sec_is0[27] &  sec_is0[28] &  sec_is0[29]
		 &  sec_is0[30]) |
		(~pri_is0[0] &  pri_is0[1] &  pri_is0[2] &  pri_is0[3]
		 &  pri_is0[4] &  pri_is0[5] &  sec_is0[21]
		 & ~sec_is0[22] &  sec_is0[26] & ~sec_is0[27]
		 &  sec_is0[28] &  sec_is0[29] &  sec_is0[30]) |
		(~pri_is0[0] &  pri_is0[1] &  pri_is0[2] &  pri_is0[3]
		 &  pri_is0[4] &  pri_is0[5] &  sec_is0[21]
		 & ~sec_is0[23] &  sec_is0[24] &  sec_is0[26]
		 & ~sec_is0[27] &  sec_is0[28] &  sec_is0[29]
		 &  sec_is0[30]) |
		(~pri_is0[0] &  pri_is0[1] &  pri_is0[2] &  pri_is0[3]
		 &  pri_is0[4] &  pri_is0[5] &  sec_is0[21]
		 & ~sec_is0[22] &  sec_is0[24] &  sec_is0[26]
		 &  sec_is0[28] &  sec_is0[29] &  sec_is0[30]) |
		( pri_is0[0] &  pri_is0[1] & ~pri_is0[2]);

assign st_is0 =  (~pri_is0[0] &  pri_is0[1] &  pri_is0[2] &  pri_is0[3]
		 &  pri_is0[4] &  pri_is0[5] &  sec_is0[20]
		 & ~sec_is0[21] & ~sec_is0[22] & ~sec_is0[23]
		 &  sec_is0[24] & ~sec_is0[26] & ~sec_is0[27]
		 & ~sec_is0[28] &  sec_is0[29] &  sec_is0[30]) |
	(~pri_is0[0] &  pri_is0[1] &  pri_is0[2] &  pri_is0[3]
	 &  pri_is0[4] &  pri_is0[5] &  sec_is0[21] & ~sec_is0[22]
	 &  sec_is0[23] &  sec_is0[24] &  sec_is0[25] &  sec_is0[26]
	 &  sec_is0[27] &  sec_is0[28] &  sec_is0[29]) |
	(~pri_is0[0] &  pri_is0[1] &  pri_is0[2] &  pri_is0[3]
	 &  pri_is0[4] &  pri_is0[5] &  sec_is0[21] & ~sec_is0[22]
	 &  sec_is0[23] &  sec_is0[24] & ~sec_is0[25] &  sec_is0[26]
	 &  sec_is0[27] &  sec_is0[28] &  sec_is0[30]) |
	(~pri_is0[0] &  pri_is0[1] &  pri_is0[2] &  pri_is0[3]
	 &  pri_is0[4] &  pri_is0[5] &  sec_is0[21] &  sec_is0[23]
	 &  sec_is0[24] & ~sec_is0[25] &  sec_is0[26] & ~sec_is0[27]
	 &  sec_is0[28] &  sec_is0[29] &  sec_is0[30]) |
	(~pri_is0[0] &  pri_is0[1] &  pri_is0[2] &  pri_is0[3]
	 &  pri_is0[4] &  pri_is0[5] &  sec_is0[21] & ~sec_is0[22]
	 &  sec_is0[23] &  sec_is0[26] & ~sec_is0[27] &  sec_is0[28]
	 &  sec_is0[29] &  sec_is0[30]) |
	( pri_is0[0] &  pri_is0[1] & ~pri_is0[2] &  pri_is0[3]);

assign indexed =  ( pri_is0[2] &  sec_is0[20] & ~sec_is0[23] & ~sec_is0[25]
	 & ~sec_is0[26] & ~sec_is0[27] & ~sec_is0[28] &  sec_is0[29]
	 &  sec_is0[30]) |
	(~pri_is0[0] &  sec_is0[21] &  sec_is0[25] &  sec_is0[26]
	 & ~sec_is0[27] &  sec_is0[28] &  sec_is0[29] &  sec_is0[30]) |
	(~pri_is0[0] &  sec_is0[21] &  sec_is0[24] &  sec_is0[26]
	 & ~sec_is0[27] &  sec_is0[28] &  sec_is0[29] &  sec_is0[30]) |
	(~pri_is0[0] &  sec_is0[21] & ~sec_is0[22] & ~sec_is0[25]
	 &  sec_is0[29]);

assign update_form =  (~pri_is0[0] &  pri_is0[1] &  pri_is0[2] &  pri_is0[3]
	 &  pri_is0[4] &  pri_is0[5] &  sec_is0[21] & ~sec_is0[22]
	 &  sec_is0[25] &  sec_is0[26] & ~sec_is0[27] &  sec_is0[28]
	 &  sec_is0[29] &  sec_is0[30]) |
		( pri_is0[0] &  pri_is0[1] & ~pri_is0[2] &  pri_is0[5]);

assign forcealign =  ( pri_is0[2] &  pri_is0[3] &  pri_is0[4] &  sec_is0[21]
		 &  sec_is0[22] &  sec_is0[23] &  sec_is0[24]
		 &  sec_is0[25] &  sec_is0[26]);

assign single_precision_ldst =  ( pri_is0[1] & ~pri_is0[2] & ~pri_is0[4]) |
		(~pri_is0[0] &  sec_is0[21] & ~sec_is0[22]
		 &  sec_is0[28] &  sec_is0[29] & ~sec_is0[30]) |
		(~pri_is0[0] &  sec_is0[21] & ~sec_is0[22]
		 & ~sec_is0[24]);

assign int_word_ldst =  ( pri_is0[2] &  sec_is0[20] & ~sec_is0[22]
		 & ~sec_is0[23] & ~sec_is0[26] & ~sec_is0[27]
		 & ~sec_is0[28] &  sec_is0[29] &  sec_is0[30]) |
		(~pri_is0[0] &  sec_is0[22] &  sec_is0[24]
		 &  sec_is0[26] & ~sec_is0[27] &  sec_is0[28]
		 &  sec_is0[29] &  sec_is0[30]) |
		(~pri_is0[0] &  sec_is0[21] & ~sec_is0[22]
		 & ~sec_is0[23] &  sec_is0[28] & ~sec_is0[29]) |
		(~pri_is0[0] &  sec_is0[21] & ~sec_is0[25]
		 & ~sec_is0[29]);

assign sign_ext_ldst =  (~pri_is0[0] &  sec_is0[21] & ~sec_is0[22]
		 & ~sec_is0[23] &  sec_is0[28] & ~sec_is0[29]
		 & ~sec_is0[30]) |
		(~pri_is0[0] &  sec_is0[22] & ~sec_is0[23]
		 &  sec_is0[24] & ~sec_is0[25]);

assign ldst_extpid =  (~pri_is0[0] &  pri_is0[1] &  pri_is0[2] &  pri_is0[3]
		 &  pri_is0[4] &  pri_is0[5] &  sec_is0[21]
		 & ~sec_is0[22] &  sec_is0[24] & ~sec_is0[25]
		 &  sec_is0[26] &  sec_is0[27] &  sec_is0[28]
		 &  sec_is0[29] &  sec_is0[30]);

assign io_port =  (~pri_is0[0] &  pri_is0[1] &  pri_is0[2] &  pri_is0[3]
		 &  pri_is0[4] &  pri_is0[5] &  sec_is0[20]
		 & ~sec_is0[21] & ~sec_is0[22] & ~sec_is0[23]
		 & ~sec_is0[26] & ~sec_is0[27] & ~sec_is0[28]
		 &  sec_is0[29] &  sec_is0[30]);

assign io_port_ext =  (~pri_is0[0] &  pri_is0[1] &  pri_is0[2] &  pri_is0[3]
		 &  pri_is0[4] &  pri_is0[5] &  sec_is0[20]
		 & ~sec_is0[21] & ~sec_is0[22] & ~sec_is0[23]
		 & ~sec_is0[25] & ~sec_is0[26] & ~sec_is0[27]
		 & ~sec_is0[28] &  sec_is0[29] &  sec_is0[30]);

assign size[0] =  (~pri_is0[1] & ~pri_is0[3]);

assign size[1] =  (~pri_is0[1] & ~pri_is0[3]);

assign size[2] =  ( pri_is0[4] &  sec_is0[21] & ~sec_is0[22] & ~sec_is0[25]
		 &  sec_is0[27] &  sec_is0[29]) |
	( pri_is0[4] &  sec_is0[21] & ~sec_is0[22] &  sec_is0[24]
	 & ~sec_is0[27]) |
	(~pri_is0[2] &  pri_is0[4]);

assign size[3] =  ( pri_is0[2] &  pri_is0[4] &  sec_is0[21] & ~sec_is0[22]
	 & ~sec_is0[24]) |
	( pri_is0[2] &  sec_is0[22] &  sec_is0[24] &  sec_is0[26]
	 & ~sec_is0[27] &  sec_is0[28] &  sec_is0[29] &  sec_is0[30]) |
	( pri_is0[1] & ~pri_is0[2] & ~pri_is0[4]);

assign size[4] =  (~pri_is0[1] & ~pri_is0[3]);

assign size[5] =  (~pri_is0[1] & ~pri_is0[3]);

assign cr_writer =  ( pri_is0[2] &  sec_is0[20] & ~sec_is0[22] & ~sec_is0[23]
	 & ~sec_is0[26] & ~sec_is0[27] & ~sec_is0[28] &  sec_is0[29]
	 &  sec_is0[30] &  sec_is0[31]) |
		( pri_is0[0] &  pri_is0[2] & ~sec_is0[25] & ~sec_is0[26]
		 & ~sec_is0[29] & ~sec_is0[30] &  sec_is0[31]) |
		( pri_is0[0] &  pri_is0[2] & ~sec_is0[21] &  sec_is0[24]
		 &  sec_is0[27] &  sec_is0[31]) |
		( pri_is0[0] &  pri_is0[2] & ~sec_is0[23] & ~sec_is0[26]
		 &  sec_is0[31]) |
		( pri_is0[0] &  pri_is0[2] &  pri_is0[4] & ~sec_is0[22]
		 & ~sec_is0[26] & ~sec_is0[27] & ~sec_is0[28]
		 & ~sec_is0[29] & ~sec_is0[30]) |
		( pri_is0[0] &  pri_is0[2] & ~sec_is0[25] &  sec_is0[28]
		 &  sec_is0[29] &  sec_is0[31]) |
		( pri_is0[2] &  sec_is0[22] & ~sec_is0[24]
		 &  sec_is0[27] &  sec_is0[31]) |
		( pri_is0[0] &  pri_is0[2] &  sec_is0[26] &  sec_is0[30]
		 &  sec_is0[31]) |
		( pri_is0[0] &  pri_is0[2] &  sec_is0[26] &  sec_is0[29]
		 &  sec_is0[31]) |
		( pri_is0[0] &  pri_is0[2] &  sec_is0[26] &  sec_is0[28]
		 &  sec_is0[31]) |
		( pri_is0[0] &  pri_is0[2] &  sec_is0[26] &  sec_is0[27]
		 &  sec_is0[31]);

assign mffgpr =  (~pri_is0[0] &  pri_is0[1] &  pri_is0[2] &  pri_is0[3]
		 &  pri_is0[4] &  pri_is0[5] &  sec_is0[20]
		 & ~sec_is0[21] & ~sec_is0[22] & ~sec_is0[23]
		 & ~sec_is0[24] & ~sec_is0[26] & ~sec_is0[27]
		 & ~sec_is0[28] &  sec_is0[29] &  sec_is0[30]) |
	(~pri_is0[0] &  pri_is0[1] &  pri_is0[2] &  pri_is0[3]
	 &  pri_is0[4] &  pri_is0[5] &  sec_is0[21] & ~sec_is0[22]
	 & ~sec_is0[23] &  sec_is0[24] &  sec_is0[25] &  sec_is0[26]
	 &  sec_is0[27] &  sec_is0[28]);

assign mftgpr =  (~pri_is0[0] &  pri_is0[1] &  pri_is0[2] &  pri_is0[3]
	 &  pri_is0[4] &  pri_is0[5] &  sec_is0[21] & ~sec_is0[22]
	 &  sec_is0[23] &  sec_is0[24] & ~sec_is0[25] &  sec_is0[26]
	 &  sec_is0[27] &  sec_is0[28] & ~sec_is0[29] &  sec_is0[30]) |
	(~pri_is0[0] &  pri_is0[1] &  pri_is0[2] &  pri_is0[3]
	 &  pri_is0[4] &  pri_is0[5] &  sec_is0[21] & ~sec_is0[22]
	 &  sec_is0[23] &  sec_is0[24] &  sec_is0[25] &  sec_is0[26]
	 &  sec_is0[27] &  sec_is0[28] &  sec_is0[29]) |
	(~pri_is0[0] &  pri_is0[1] &  pri_is0[2] &  pri_is0[3]
	 &  pri_is0[4] &  pri_is0[5] &  sec_is0[20] & ~sec_is0[21]
	 & ~sec_is0[22] & ~sec_is0[23] &  sec_is0[24] & ~sec_is0[26]
	 & ~sec_is0[27] & ~sec_is0[28] &  sec_is0[29] &  sec_is0[30]);

assign fdiv_is0 =  ( pri_is0[0] &  pri_is0[1] &  pri_is0[2] &  pri_is0[4]
	 &  pri_is0[5] &  sec_is0[26] & ~sec_is0[27] & ~sec_is0[28]
	 &  sec_is0[29] & ~sec_is0[30]);

assign fsqrt_is0 =  ( pri_is0[0] &  pri_is0[1] &  pri_is0[2] &  pri_is0[4]
	 &  pri_is0[5] &  sec_is0[26] & ~sec_is0[27] &  sec_is0[28]
	 &  sec_is0[29] & ~sec_is0[30]);

assign only_from_ucode =  (~pri_is0[0] &  pri_is0[1] &  pri_is0[2] &  pri_is0[3]
	 &  pri_is0[4] &  pri_is0[5] &  sec_is0[21] & ~sec_is0[22]
	 &  sec_is0[24] &  sec_is0[25] &  sec_is0[26] &  sec_is0[27]
	 &  sec_is0[28] &  sec_is0[29]) |
		(~pri_is0[0] &  pri_is0[1] &  pri_is0[2] &  pri_is0[3]
		 &  pri_is0[4] &  pri_is0[5] &  sec_is0[21]
		 & ~sec_is0[22] &  sec_is0[23] &  sec_is0[24]
		 & ~sec_is0[25] &  sec_is0[26] &  sec_is0[27]
		 &  sec_is0[28] & ~sec_is0[29] &  sec_is0[30]) |
		(~pri_is0[0] &  pri_is0[1] &  pri_is0[2] &  pri_is0[3]
		 &  pri_is0[4] &  pri_is0[5] &  sec_is0[21]
		 & ~sec_is0[22] & ~sec_is0[23] &  sec_is0[24]
		 &  sec_is0[25] &  sec_is0[26] &  sec_is0[27]
		 &  sec_is0[28]) |
		( pri_is0[0] &  pri_is0[1] &  pri_is0[2] &  pri_is0[4]
		 &  pri_is0[5] &  sec_is0[26] & ~sec_is0[27]
		 & ~sec_is0[28] & ~sec_is0[29] &  sec_is0[30]) |
		( pri_is0[0] &  pri_is0[1] &  pri_is0[2] &  pri_is0[3]
		 &  pri_is0[4] &  pri_is0[5] &  sec_is0[26]
		 & ~sec_is0[27] & ~sec_is0[28] & ~sec_is0[29]);

assign no_ram =  (~pri_is0[0] &  pri_is0[1] &  pri_is0[2] &  pri_is0[3]
		 &  pri_is0[4] &  pri_is0[5] &  sec_is0[21]
		 & ~sec_is0[22] & ~sec_is0[23] &  sec_is0[25]
		 &  sec_is0[26] & ~sec_is0[27] &  sec_is0[28]
		 &  sec_is0[29] &  sec_is0[30]) |
	( pri_is0[0] &  pri_is0[1] & ~pri_is0[2] & ~pri_is0[3]
	 &  pri_is0[5]);

assign only_graphics_mode =  ( pri_is0[0] &  pri_is0[1] &  pri_is0[2]
	 & ~pri_is0[3] &  pri_is0[4] &  pri_is0[5] & ~sec_is0[21]
	 & ~sec_is0[22] &  sec_is0[23] &  sec_is0[24] & ~sec_is0[26]
	 & ~sec_is0[27] &  sec_is0[28] & ~sec_is0[29] &  sec_is0[30]
	 & ~sec_is0[31]) |
		(~pri_is0[0] &  pri_is0[1] &  pri_is0[2] &  pri_is0[3]
		 &  pri_is0[4] &  pri_is0[5] &  sec_is0[21]
		 & ~sec_is0[22] & ~sec_is0[23] &  sec_is0[24]
		 &  sec_is0[25] &  sec_is0[26] &  sec_is0[27]
		 &  sec_is0[28]) |
		(~pri_is0[0] &  pri_is0[1] &  pri_is0[2] &  pri_is0[3]
		 &  pri_is0[4] &  pri_is0[5] &  sec_is0[21]
		 & ~sec_is0[22] &  sec_is0[23] &  sec_is0[24]
		 & ~sec_is0[25] &  sec_is0[26] &  sec_is0[27]
		 &  sec_is0[28] & ~sec_is0[29] &  sec_is0[30]) |
		(~pri_is0[0] &  pri_is0[1] &  pri_is0[2] &  pri_is0[3]
		 &  pri_is0[4] &  pri_is0[5] &  sec_is0[21]
		 & ~sec_is0[22] &  sec_is0[24] &  sec_is0[25]
		 &  sec_is0[26] &  sec_is0[27] &  sec_is0[28]
		 &  sec_is0[29]);

//@@ ESPRESSO LOGIC END @@



      assign ldst_tag = {single_precision_ldst, int_word_ldst, sign_ext_ldst, iu_au_iu4_ucode_ext[0], ldst_tag_addr[0:4]};		// for lfiwax

      assign ldst_tag_addr = (mftgpr == 1'b0) ? is0_instr[06:10] :
                             is0_instr[16:20];

      assign ram_mode_v = iu_au_iu4_isram;

      //----------------------------------------------------------------------------------------------------------------------
      // config bits
      assign iu_au_config_iucr_din = iu_au_config_iucr;

      assign config_reg_scin = 0;


      tri_rlmreg_p #(.INIT(0), .WIDTH(8)) config_reg(
         .vd(vdd),
         .gd(gnd),
         .force_t(force_t),
         .delay_lclkr(delay_lclkr),
         .nclk(nclk),
         .mpw1_b(mpw1_b),
         .act(tiup),
         .mpw2_b(mpw2_b),
         .thold_b(pc_iu_func_sl_thold_0_b),
         .sg(pc_iu_sg_0),
	 .d_mode(tiup),
         .scin(config_reg_scin[0:7]),
         .scout(config_reg_scout[0:7]),
         .din(iu_au_config_iucr_din),
         .dout(iu_au_config_iucr_l2)
      );

      assign iu_au_config_iucr_int[0:7] = iu_au_config_iucr_l2[0:7];

      assign graphics_mode = iu_au_config_iucr_int[0];

      assign spare_unused[4:7] = iu_au_config_iucr_int[4:7];

      assign is0_is_ucode = iu_au_iu4_ucode[0];

      assign in_ucode_mode = iu_au_iu4_ucode[0] & is0_instr_v;

      // special ucode instructions getting issued when not doing ucode is bad
      assign is0_invalid_kill_uc = ((~(in_ucode_mode | ram_mode_v)) & only_from_ucode) | ((~(graphics_mode | in_ucode_mode | ram_mode_v)) & only_graphics_mode);		// can use any graphics mode insr in ucode

      // the XU must now do something like:

      //au_iu_is0_i_dec_internal <=  (not au_iu_is0_i_dec_b) and not (not in_ucode_mode and au_iu_is0_ucode_only);

      assign is0_invalid_kill = ((~(graphics_mode | in_ucode_mode)) & only_graphics_mode) | is0_invalid_kill_uc;		// can use any graphics mode insr in ucode
      //is0_invalid_kill <=  '0';

      assign au_iu_iu4_no_ram = no_ram;

      assign is0_kill_or_divsqrt_b = (~(is0_invalid_kill));

      assign is0_i_dec_b = (~(isfu_dec_is0 & is0_kill_or_divsqrt_b));		// inverted for timing
      assign au_iu_iu4_i_dec_b = is0_i_dec_b;

      assign au_iu_is0_i_dec = (~is0_i_dec_b);
      assign spare_unused[3] = au_iu_is0_i_dec;

      // fdiv and fsqrt will be handled by ucode.  The fu may issue them lateer
      // This signal is passed down the pipe to rf1, because
      // these opcodes are used to initiate some operand checking so they should continue down the pipe and not be flushed because of ucode.

      // During fdiv/fsqrt the axu may select this thread before or after the "real" fxu selection.
      // If the axu selects this thread earlier than the fxu, s1 is simply updated early.
      // If the axu selects this thread later than the fxu, ucode instructions would get wiped out by the flush
      // This signal protects the instruction from being flushed
      //ignore_flush_is0 <= (fdiv_is0 or fsqrt_is0) and isfu_dec_is0;  -- these opcodes will not change the FpScr or any Fpr.  Only scratch reg s0 will be changed
      assign ignore_flush_is0 = 1'b0;		// disabled for a2o

      //----------------------------------------------------------------------------------------------------------------------

      assign is0_to_ucode = (iu_au_iu4_2ucode) & isfu_dec_is0;		//uCode from either a denorm or fdiv(s)(.) or fsqrt(s)(.)
      assign au_iu_iu4_ucode[0:2] = iu_au_iu4_ucode[0:2];

      assign is0_ldst_ra = (mftgpr == 1'b0) ? {iu_au_iu4_ucode_ext[1], is0_instr[11:15]} :
                           {iu_au_iu4_ucode_ext[0], is0_instr[6:10]};		// for mftgpr, make RA the target, same as updates

      assign is0_zero_r0 = ld_st_is0 & (is0_ldst_ra == 6'b000000);

      //----------------------------------------------------------------------------------------------------------------------
      // Interface to Core Decode

      // mftgpr RT,   FRB
      //        6:10, 16:20
      // mffgpr FRT,  RB
      //        6:10, 16:20
      // mfdp   FRT     t2     (mffgpr and io_port)
      //        6:10
      // mtdp   FRS     s3     (mftgpr and io_port)
      //        6:10
      // lfdx   FRT, RA,RB
      //        6:10,11:15,16:20
      // stfdx  FRS, RA,RB
      //        6:10,11:15,16:20

      assign au_iu_iu4_t1_v = (update_form | mftgpr | fpscr_wr) & (~iu_au_iu4_ucode[1]);
      assign au_iu_iu4_t1_t[0:2] = (fpscr_wr == 1'b1) ? 3'b111 : 		//fpscr or gpr
                                   3'b000;
      assign au_iu_iu4_t1_a6[0:5] = (({iu_au_iu4_ucode_ext[1], is0_instr[11:15]}) & ({6{(~mftgpr) & (~fpscr_wr)}})) |
                                    (({iu_au_iu4_ucode_ext[0], is0_instr[6:10]})  & ({6{  mftgpr  & (~fpscr_wr)}})) |
	                            ((6'b000000) & ({6{fpscr_wr}}));

      //----------------------------------------------------------------------------------------------------------------------
      assign au_iu_iu4_t2_v = tv & (~iu_au_iu4_ucode[1]);
      assign au_iu_iu4_t2_a6[0:5] = (tv == 1'b0 & fpscr_wr == 1'b1) ? 6'b110000 : 		//for compares, need fpscr rename, big targ
                                    {iu_au_iu4_ucode_ext[0], is0_instr[06:10]};
      assign au_iu_iu4_t2_t[0:2] = 3'b110;		//fpr

      //----------------------------------------------------------------------------------------------------------------------
      assign au_iu_iu4_t3_v = cr_writer & (~iu_au_iu4_ucode[1]);
      assign au_iu_iu4_t3_a6[0:5] = ({3'b000, is0_instr[06:08]} & {6{(~record_form)}}) | ((6'b000001) & {6{record_form}});
      assign au_iu_iu4_t3_t[0:2] = 3'b001;		//cr

      //----------------------------------------------------------------------------------------------------------------------
      assign au_iu_iu4_s1_v = ((ld_st_is0 & (~is0_zero_r0) & (~mftgpr) & (~mffgpr)) & ld_st_is0) | (av & (~ld_st_is0));
      assign au_iu_iu4_s1_a6[0:5] = ((is0_ldst_ra[0:5]) & {6{ld_st_is0}}) | (({iu_au_iu4_ucode_ext[1], is0_instr[11:15]}) & {6{(~ld_st_is0)}});

      //gpr
	assign au_iu_iu4_s1_t[0:2] = (3'b000 & {3{ld_st_is0}}) | (3'b110 & {3{(~ld_st_is0)}});		//fpr

      //----------------------------------------------------------------------------------------------------------------------
      assign au_iu_iu4_s2_v = ((indexed | mffgpr) & ld_st_is0) | (bv & (~ld_st_is0));
      assign au_iu_iu4_s2_a6[0:5] = {iu_au_iu4_ucode_ext[2], is0_instr[16:20]};
      //gpr
	assign au_iu_iu4_s2_t[0:2] = (3'b000 & {3{ld_st_is0}}) | (3'b110 & {3{(~ld_st_is0)}});		//fpr

      //----------------------------------------------------------------------------------------------------------------------
      assign au_iu_iu4_s3_v = (st_is0 & (~mftgpr) & ld_st_is0) | (cv & (~ld_st_is0));
	assign au_iu_iu4_s3_a6[0:5] = (({iu_au_iu4_ucode_ext[0], is0_instr[06:10]}) & {6{ld_st_is0 & (~(mffgpr | mftgpr))}}) |
	                              (({iu_au_iu4_ucode_ext[2], is0_instr[16:20]}) & {6{ld_st_is0 & (  mffgpr | mftgpr) }}) |
	                              (({iu_au_iu4_ucode_ext[3], is0_instr[21:25]}) & {6{(~ld_st_is0)}});
      //gpr
	assign au_iu_iu4_s3_t[0:2] = (3'b000 & {3{mffgpr}}) | (3'b110 & {3{(~mffgpr)}});		//fpr

      //----------------------------------------------------------------------------------------------------------------------
      generate
         if (`GPR_POOL_ENC > 6)
         begin : gpr_pool
            assign au_iu_iu4_t1_a[0:`GPR_POOL_ENC - 7] = 0;
            assign au_iu_iu4_t2_a[0:`GPR_POOL_ENC - 7] = 0;
            assign au_iu_iu4_t3_a[0:`GPR_POOL_ENC - 7] = 0;
            assign au_iu_iu4_s1_a[0:`GPR_POOL_ENC - 7] = 0;
            assign au_iu_iu4_s2_a[0:`GPR_POOL_ENC - 7] = 0;
            assign au_iu_iu4_s3_a[0:`GPR_POOL_ENC - 7] = 0;
         end
      endgenerate
      assign au_iu_iu4_t1_a[`GPR_POOL_ENC - 6:`GPR_POOL_ENC - 1] = au_iu_iu4_t1_a6[0:5];
      assign au_iu_iu4_t2_a[`GPR_POOL_ENC - 6:`GPR_POOL_ENC - 1] = au_iu_iu4_t2_a6[0:5];
      assign au_iu_iu4_t3_a[`GPR_POOL_ENC - 6:`GPR_POOL_ENC - 1] = au_iu_iu4_t3_a6[0:5];
      assign au_iu_iu4_s1_a[`GPR_POOL_ENC - 6:`GPR_POOL_ENC - 1] = au_iu_iu4_s1_a6[0:5];
      assign au_iu_iu4_s2_a[`GPR_POOL_ENC - 6:`GPR_POOL_ENC - 1] = au_iu_iu4_s2_a6[0:5];
      assign au_iu_iu4_s3_a[`GPR_POOL_ENC - 6:`GPR_POOL_ENC - 1] = au_iu_iu4_s3_a6[0:5];

      //----------------------------------------------------------------------------------------------------------------------
      assign isLoad = ld_st_is0 & (~st_is0) & (~(mffgpr | mftgpr));
      assign isStore = ld_st_is0 & (st_is0 | mftgpr) & (~mffgpr);

      assign au_iu_iu4_isload = isLoad;
      assign au_iu_iu4_isstore = isStore;

      assign au_iu_iu4_ilat[0:2] = (3'b100 & {3{ld_st_is0 & (~st_is0)}}) | (3'b011 & {3{ld_st_is0 & st_is0 & (~mftgpr)}}) | (3'b110 & {3{ld_st_is0 & st_is0 & mftgpr}}) | (3'b110 & {3{(~ld_st_is0)}});
      assign au_iu_iu4_ord = ordered & (~iu_au_iu4_ucode[1]);
      assign au_iu_iu4_cord = cordered & (~iu_au_iu4_ucode[1]);

      assign au_iu_iu4_spec = ld_st_is0;

      // To set the ESR bits
      assign au_iu_iu4_type_fp = isfu_dec_is0;
      assign au_iu_iu4_type_ap = 1'b0;
      assign au_iu_iu4_type_spv = 1'b0;
      assign au_iu_iu4_type_st = st_is0;

      assign au_iu_iu4_rte_lq = ld_st_is0;
      assign au_iu_iu4_rte_sq = isStore;
      assign au_iu_iu4_rte_axu0 = isfu_dec_is0 & (~(ld_st_is0 & (~st_is0))) & ~(isStore & iu_au_iu4_ucode[1]); //don't route to axu on a store pressissue
      assign au_iu_iu4_rte_axu1 = 1'b0;

      assign au_iu_iu4_async_block = fpscr_mv;

      //----------------------------------------------------------------------------------------------------------------------

      assign i_dec_so = 1'b0;
      assign fu_dec_debug = 0;


endmodule
