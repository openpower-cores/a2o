// © IBM Corp. 2020
// This softcore is licensed under and subject to the terms of the CC-BY 4.0
// license (https://creativecommons.org/licenses/by/4.0/legalcode). 
// Additional rights, including the right to physically implement a softcore 
// that is compliant with the required sections of the Power ISA 
// Specification, will be available at no cost via the OpenPOWER Foundation. 
// This README will be updated with additional information when OpenPOWER's 
// license is available.

`timescale 1 ns / 1 ns

//  Description:  Completion Unit
//
//*****************************************************************************

`include "tri_a2o.vh"

module iuq_cpl_top(
   // Clocks
    (* pin_data="PIN_FUNCTION=/G_CLK/" *)
   input [0:`NCLK_WIDTH-1]    nclk,

   // Pervasive
   input                       tc_ac_ccflush_dc,
   input                       clkoff_dc_b,
   input                       d_mode_dc,
   input                       delay_lclkr_dc,
   input                       mpw1_dc_b,
   input                       mpw2_dc_b,
   input                       pc_iu_func_sl_thold_2,
   input                       pc_iu_func_slp_sl_thold_2,
   input                       pc_iu_sg_2,
   input [0:`THREADS]          cp_scan_in,
   output [0:`THREADS]         cp_scan_out,

   // Perfomance selectors
   input                       pc_iu_event_bus_enable,
   input [0:2]		       pc_iu_event_count_mode,

   input [0:31]                spr_cp_perf_event_mux_ctrls,
   input [0:4*`THREADS-1]      event_bus_in,
   output [0:4*`THREADS-1]     event_bus_out,

   // Instruction 0 Issue
   input                       rn_cp_iu6_t0_i0_vld,
   input [1:`ITAG_SIZE_ENC-1]  rn_cp_iu6_t0_i0_itag,
   input [0:2]                 rn_cp_iu6_t0_i0_ucode,
   input                       rn_cp_iu6_t0_i0_fuse_nop,
   input                       rn_cp_iu6_t0_i0_rte_lq,
   input                       rn_cp_iu6_t0_i0_rte_sq,
   input                       rn_cp_iu6_t0_i0_rte_fx0,
   input                       rn_cp_iu6_t0_i0_rte_fx1,
   input                       rn_cp_iu6_t0_i0_rte_axu0,
   input                       rn_cp_iu6_t0_i0_rte_axu1,

   input [62-`EFF_IFAR_WIDTH:61] rn_cp_iu6_t0_i0_ifar,
   input [62-`EFF_IFAR_WIDTH:61] rn_cp_iu6_t0_i0_bta,
   input                       rn_cp_iu6_t0_i0_isram,
   input [0:31]                rn_cp_iu6_t0_i0_instr,

   input                       rn_cp_iu6_t0_i0_valop,
   input [0:2]                 rn_cp_iu6_t0_i0_error,
   input                       rn_cp_iu6_t0_i0_br_pred,
   input                       rn_cp_iu6_t0_i0_bh_update,
   input [0:1]                 rn_cp_iu6_t0_i0_bh0_hist,
   input [0:1]                 rn_cp_iu6_t0_i0_bh1_hist,
   input [0:1]                 rn_cp_iu6_t0_i0_bh2_hist,
   input [0:9]                 rn_cp_iu6_t0_i0_gshare,
   input [0:2]                 rn_cp_iu6_t0_i0_ls_ptr,
   input                       rn_cp_iu6_t0_i0_match,

   input                       rn_cp_iu6_t0_i0_type_fp,
   input                       rn_cp_iu6_t0_i0_type_ap,
   input                       rn_cp_iu6_t0_i0_type_spv,
   input                       rn_cp_iu6_t0_i0_type_st,
   input                       rn_cp_iu6_t0_i0_async_block,
   input                       rn_cp_iu6_t0_i0_np1_flush,

   input                       rn_cp_iu6_t0_i0_t1_v,
   input [0:2]                 rn_cp_iu6_t0_i0_t1_t,
   input [0:`GPR_POOL_ENC-1]   rn_cp_iu6_t0_i0_t1_p,
   input [0:`GPR_POOL_ENC-1]   rn_cp_iu6_t0_i0_t1_a,

   input                       rn_cp_iu6_t0_i0_t2_v,
   input [0:2]                 rn_cp_iu6_t0_i0_t2_t,
   input [0:`GPR_POOL_ENC-1]   rn_cp_iu6_t0_i0_t2_p,
   input [0:`GPR_POOL_ENC-1]   rn_cp_iu6_t0_i0_t2_a,

   input                       rn_cp_iu6_t0_i0_t3_v,
   input [0:2]                 rn_cp_iu6_t0_i0_t3_t,
   input [0:`GPR_POOL_ENC-1]   rn_cp_iu6_t0_i0_t3_p,
   input [0:`GPR_POOL_ENC-1]   rn_cp_iu6_t0_i0_t3_a,

   input                       rn_cp_iu6_t0_i0_btb_entry,
   input [0:1]                 rn_cp_iu6_t0_i0_btb_hist,
   input                       rn_cp_iu6_t0_i0_bta_val,

   // Instruction 1 Issue
   input                       rn_cp_iu6_t0_i1_vld,
   input [1:`ITAG_SIZE_ENC-1]  rn_cp_iu6_t0_i1_itag,
   input [0:2]                 rn_cp_iu6_t0_i1_ucode,
   input                       rn_cp_iu6_t0_i1_fuse_nop,
   input                       rn_cp_iu6_t0_i1_rte_lq,
   input                       rn_cp_iu6_t0_i1_rte_sq,
   input                       rn_cp_iu6_t0_i1_rte_fx0,
   input                       rn_cp_iu6_t0_i1_rte_fx1,
   input                       rn_cp_iu6_t0_i1_rte_axu0,
   input                       rn_cp_iu6_t0_i1_rte_axu1,

   input [62-`EFF_IFAR_WIDTH:61] rn_cp_iu6_t0_i1_ifar,
   input [62-`EFF_IFAR_WIDTH:61] rn_cp_iu6_t0_i1_bta,
   input                       rn_cp_iu6_t0_i1_isram,
   input [0:31]                rn_cp_iu6_t0_i1_instr,

   input                       rn_cp_iu6_t0_i1_valop,
   input [0:2]                 rn_cp_iu6_t0_i1_error,
   input                       rn_cp_iu6_t0_i1_br_pred,
   input                       rn_cp_iu6_t0_i1_bh_update,
   input [0:1]                 rn_cp_iu6_t0_i1_bh0_hist,
   input [0:1]                 rn_cp_iu6_t0_i1_bh1_hist,
   input [0:1]                 rn_cp_iu6_t0_i1_bh2_hist,
   input [0:9]                 rn_cp_iu6_t0_i1_gshare,
   input [0:2]                 rn_cp_iu6_t0_i1_ls_ptr,
   input                       rn_cp_iu6_t0_i1_match,

   input                       rn_cp_iu6_t0_i1_type_fp,
   input                       rn_cp_iu6_t0_i1_type_ap,
   input                       rn_cp_iu6_t0_i1_type_spv,
   input                       rn_cp_iu6_t0_i1_type_st,
   input                       rn_cp_iu6_t0_i1_async_block,
   input                       rn_cp_iu6_t0_i1_np1_flush,

   input                       rn_cp_iu6_t0_i1_t1_v,
   input [0:2]                 rn_cp_iu6_t0_i1_t1_t,
   input [0:`GPR_POOL_ENC-1]   rn_cp_iu6_t0_i1_t1_p,
   input [0:`GPR_POOL_ENC-1]   rn_cp_iu6_t0_i1_t1_a,

   input                       rn_cp_iu6_t0_i1_t2_v,
   input [0:2]                 rn_cp_iu6_t0_i1_t2_t,
   input [0:`GPR_POOL_ENC-1]   rn_cp_iu6_t0_i1_t2_p,
   input [0:`GPR_POOL_ENC-1]   rn_cp_iu6_t0_i1_t2_a,

   input                       rn_cp_iu6_t0_i1_t3_v,
   input [0:2]                 rn_cp_iu6_t0_i1_t3_t,
   input [0:`GPR_POOL_ENC-1]   rn_cp_iu6_t0_i1_t3_p,
   input [0:`GPR_POOL_ENC-1]   rn_cp_iu6_t0_i1_t3_a,

   input                       rn_cp_iu6_t0_i1_btb_entry,
   input [0:1]                 rn_cp_iu6_t0_i1_btb_hist,
   input                       rn_cp_iu6_t0_i1_bta_val,

`ifndef THREADS1
   // Instruction 0 Issue
   input                       rn_cp_iu6_t1_i0_vld,
   input [1:`ITAG_SIZE_ENC-1]  rn_cp_iu6_t1_i0_itag,
   input [0:2]                 rn_cp_iu6_t1_i0_ucode,
   input                       rn_cp_iu6_t1_i0_fuse_nop,
   input                       rn_cp_iu6_t1_i0_rte_lq,
   input                       rn_cp_iu6_t1_i0_rte_sq,
   input                       rn_cp_iu6_t1_i0_rte_fx0,
   input                       rn_cp_iu6_t1_i0_rte_fx1,
   input                       rn_cp_iu6_t1_i0_rte_axu0,
   input                       rn_cp_iu6_t1_i0_rte_axu1,

   input [62-`EFF_IFAR_WIDTH:61] rn_cp_iu6_t1_i0_ifar,
   input [62-`EFF_IFAR_WIDTH:61] rn_cp_iu6_t1_i0_bta,
   input                       rn_cp_iu6_t1_i0_isram,
   input [0:31]                rn_cp_iu6_t1_i0_instr,

   input                       rn_cp_iu6_t1_i0_valop,
   input [0:2]                 rn_cp_iu6_t1_i0_error,
   input                       rn_cp_iu6_t1_i0_br_pred,
   input                       rn_cp_iu6_t1_i0_bh_update,
   input [0:1]                 rn_cp_iu6_t1_i0_bh0_hist,
   input [0:1]                 rn_cp_iu6_t1_i0_bh1_hist,
   input [0:1]                 rn_cp_iu6_t1_i0_bh2_hist,
   input [0:9]                 rn_cp_iu6_t1_i0_gshare,
   input [0:2]                 rn_cp_iu6_t1_i0_ls_ptr,
   input                       rn_cp_iu6_t1_i0_match,

   input                       rn_cp_iu6_t1_i0_type_fp,
   input                       rn_cp_iu6_t1_i0_type_ap,
   input                       rn_cp_iu6_t1_i0_type_spv,
   input                       rn_cp_iu6_t1_i0_type_st,
   input                       rn_cp_iu6_t1_i0_async_block,
   input                       rn_cp_iu6_t1_i0_np1_flush,

   input                       rn_cp_iu6_t1_i0_t1_v,
   input [0:2]                 rn_cp_iu6_t1_i0_t1_t,
   input [0:`GPR_POOL_ENC-1]   rn_cp_iu6_t1_i0_t1_p,
   input [0:`GPR_POOL_ENC-1]   rn_cp_iu6_t1_i0_t1_a,

   input                       rn_cp_iu6_t1_i0_t2_v,
   input [0:2]                 rn_cp_iu6_t1_i0_t2_t,
   input [0:`GPR_POOL_ENC-1]   rn_cp_iu6_t1_i0_t2_p,
   input [0:`GPR_POOL_ENC-1]   rn_cp_iu6_t1_i0_t2_a,

   input                       rn_cp_iu6_t1_i0_t3_v,
   input [0:2]                 rn_cp_iu6_t1_i0_t3_t,
   input [0:`GPR_POOL_ENC-1]   rn_cp_iu6_t1_i0_t3_p,
   input [0:`GPR_POOL_ENC-1]   rn_cp_iu6_t1_i0_t3_a,

   input                       rn_cp_iu6_t1_i0_btb_entry,
   input [0:1]                 rn_cp_iu6_t1_i0_btb_hist,
   input                       rn_cp_iu6_t1_i0_bta_val,

   // Instruction 1 Issue
   input                       rn_cp_iu6_t1_i1_vld,
   input [1:`ITAG_SIZE_ENC-1]  rn_cp_iu6_t1_i1_itag,
   input [0:2]                 rn_cp_iu6_t1_i1_ucode,
   input                       rn_cp_iu6_t1_i1_fuse_nop,
   input                       rn_cp_iu6_t1_i1_rte_lq,
   input                       rn_cp_iu6_t1_i1_rte_sq,
   input                       rn_cp_iu6_t1_i1_rte_fx0,
   input                       rn_cp_iu6_t1_i1_rte_fx1,
   input                       rn_cp_iu6_t1_i1_rte_axu0,
   input                       rn_cp_iu6_t1_i1_rte_axu1,

   input [62-`EFF_IFAR_WIDTH:61] rn_cp_iu6_t1_i1_ifar,
   input [62-`EFF_IFAR_WIDTH:61] rn_cp_iu6_t1_i1_bta,
   input                       rn_cp_iu6_t1_i1_isram,
   input [0:31]                rn_cp_iu6_t1_i1_instr,

   input                       rn_cp_iu6_t1_i1_valop,
   input [0:2]                 rn_cp_iu6_t1_i1_error,
   input                       rn_cp_iu6_t1_i1_br_pred,
   input                       rn_cp_iu6_t1_i1_bh_update,
   input [0:1]                 rn_cp_iu6_t1_i1_bh0_hist,
   input [0:1]                 rn_cp_iu6_t1_i1_bh1_hist,
   input [0:1]                 rn_cp_iu6_t1_i1_bh2_hist,
   input [0:9]                 rn_cp_iu6_t1_i1_gshare,
   input [0:2]                 rn_cp_iu6_t1_i1_ls_ptr,
   input                       rn_cp_iu6_t1_i1_match,

   input                       rn_cp_iu6_t1_i1_type_fp,
   input                       rn_cp_iu6_t1_i1_type_ap,
   input                       rn_cp_iu6_t1_i1_type_spv,
   input                       rn_cp_iu6_t1_i1_type_st,
   input                       rn_cp_iu6_t1_i1_async_block,
   input                       rn_cp_iu6_t1_i1_np1_flush,

   input                       rn_cp_iu6_t1_i1_t1_v,
   input [0:2]                 rn_cp_iu6_t1_i1_t1_t,
   input [0:`GPR_POOL_ENC-1]   rn_cp_iu6_t1_i1_t1_p,
   input [0:`GPR_POOL_ENC-1]   rn_cp_iu6_t1_i1_t1_a,

   input                       rn_cp_iu6_t1_i1_t2_v,
   input [0:2]                 rn_cp_iu6_t1_i1_t2_t,
   input [0:`GPR_POOL_ENC-1]   rn_cp_iu6_t1_i1_t2_p,
   input [0:`GPR_POOL_ENC-1]   rn_cp_iu6_t1_i1_t2_a,

   input                       rn_cp_iu6_t1_i1_t3_v,
   input [0:2]                 rn_cp_iu6_t1_i1_t3_t,
   input [0:`GPR_POOL_ENC-1]   rn_cp_iu6_t1_i1_t3_p,
   input [0:`GPR_POOL_ENC-1]   rn_cp_iu6_t1_i1_t3_a,

   input                       rn_cp_iu6_t1_i1_btb_entry,
   input [0:1]                 rn_cp_iu6_t1_i1_btb_hist,
   input                       rn_cp_iu6_t1_i1_bta_val,
 `endif

   // completion empty
   output [0:`THREADS-1]       cp_rn_empty,
   output [0:`THREADS-1]       cp_async_block,

   // Instruction 0 Complete
   output                      cp_rn_t0_i0_v,
   output                      cp_rn_t0_i0_axu_exception_val,
   output [0:3]                cp_rn_t0_i0_axu_exception,
   output                      cp_rn_t0_i0_t1_v,
   output [0:2]                cp_rn_t0_i0_t1_t,
   output [0:`GPR_POOL_ENC-1]  cp_rn_t0_i0_t1_p,
   output [0:`GPR_POOL_ENC-1]  cp_rn_t0_i0_t1_a,

   output                      cp_rn_t0_i0_t2_v,
   output [0:2]                cp_rn_t0_i0_t2_t,
   output [0:`GPR_POOL_ENC-1]  cp_rn_t0_i0_t2_p,
   output [0:`GPR_POOL_ENC-1]  cp_rn_t0_i0_t2_a,

   output                      cp_rn_t0_i0_t3_v,
   output [0:2]                cp_rn_t0_i0_t3_t,
   output [0:`GPR_POOL_ENC-1]  cp_rn_t0_i0_t3_p,
   output [0:`GPR_POOL_ENC-1]  cp_rn_t0_i0_t3_a,

   // Instruction 1 Complete
   output                      cp_rn_t0_i1_v,
   output                      cp_rn_t0_i1_axu_exception_val,
   output [0:3]                cp_rn_t0_i1_axu_exception,
   output                      cp_rn_t0_i1_t1_v,
   output [0:2]                cp_rn_t0_i1_t1_t,
   output [0:`GPR_POOL_ENC-1]  cp_rn_t0_i1_t1_p,
   output [0:`GPR_POOL_ENC-1]  cp_rn_t0_i1_t1_a,

   output                      cp_rn_t0_i1_t2_v,
   output [0:2]                cp_rn_t0_i1_t2_t,
   output [0:`GPR_POOL_ENC-1]  cp_rn_t0_i1_t2_p,
   output [0:`GPR_POOL_ENC-1]  cp_rn_t0_i1_t2_a,

   output                      cp_rn_t0_i1_t3_v,
   output [0:2]                cp_rn_t0_i1_t3_t,
   output [0:`GPR_POOL_ENC-1]  cp_rn_t0_i1_t3_p,
   output [0:`GPR_POOL_ENC-1]  cp_rn_t0_i1_t3_a,

`ifndef THREADS1
   // Instruction 0 Complete
   output                      cp_rn_t1_i0_v,
   output                      cp_rn_t1_i0_axu_exception_val,
   output [0:3]                cp_rn_t1_i0_axu_exception,
   output                      cp_rn_t1_i0_t1_v,
   output [0:2]                cp_rn_t1_i0_t1_t,
   output [0:`GPR_POOL_ENC-1]  cp_rn_t1_i0_t1_p,
   output [0:`GPR_POOL_ENC-1]  cp_rn_t1_i0_t1_a,

   output                      cp_rn_t1_i0_t2_v,
   output [0:2]                cp_rn_t1_i0_t2_t,
   output [0:`GPR_POOL_ENC-1]  cp_rn_t1_i0_t2_p,
   output [0:`GPR_POOL_ENC-1]  cp_rn_t1_i0_t2_a,

   output                      cp_rn_t1_i0_t3_v,
   output [0:2]                cp_rn_t1_i0_t3_t,
   output [0:`GPR_POOL_ENC-1]  cp_rn_t1_i0_t3_p,
   output [0:`GPR_POOL_ENC-1]  cp_rn_t1_i0_t3_a,

   // Instruction 1 Complete
   output                      cp_rn_t1_i1_v,
   output                      cp_rn_t1_i1_axu_exception_val,
   output [0:3]                cp_rn_t1_i1_axu_exception,
   output                      cp_rn_t1_i1_t1_v,
   output [0:2]                cp_rn_t1_i1_t1_t,
   output [0:`GPR_POOL_ENC-1]  cp_rn_t1_i1_t1_p,
   output [0:`GPR_POOL_ENC-1]  cp_rn_t1_i1_t1_a,

   output                      cp_rn_t1_i1_t2_v,
   output [0:2]                cp_rn_t1_i1_t2_t,
   output [0:`GPR_POOL_ENC-1]  cp_rn_t1_i1_t2_p,
   output [0:`GPR_POOL_ENC-1]  cp_rn_t1_i1_t2_a,

   output                      cp_rn_t1_i1_t3_v,
   output [0:2]                cp_rn_t1_i1_t3_t,
   output [0:`GPR_POOL_ENC-1]  cp_rn_t1_i1_t3_p,
   output [0:`GPR_POOL_ENC-1]  cp_rn_t1_i1_t3_a,
`endif

   // Branch Prediction Complete
   output                      cp_bp_t0_val,
   output [62-`EFF_IFAR_WIDTH:61] cp_bp_t0_ifar,
   output [0:1]                cp_bp_t0_bh0_hist,
   output [0:1]                cp_bp_t0_bh1_hist,
   output [0:1]                cp_bp_t0_bh2_hist,
   output                      cp_bp_t0_br_pred,
   output                      cp_bp_t0_br_taken,
   output                      cp_bp_t0_bh_update,
   output                      cp_bp_t0_bcctr,
   output                      cp_bp_t0_bclr,
   output                      cp_bp_t0_getnia,
   output                      cp_bp_t0_group,
   output                      cp_bp_t0_lk,
   output [0:1]                cp_bp_t0_bh,
   output [0:9]                cp_bp_t0_gshare,
   output [0:2]                cp_bp_t0_ls_ptr,
   output [62-`EFF_IFAR_WIDTH:61] cp_bp_t0_ctr,
   output                      cp_bp_t0_btb_entry,
   output [0:1]                cp_bp_t0_btb_hist,

`ifndef THREADS1
   // Branch Prediction Complete
   output                      cp_bp_t1_val,
   output [62-`EFF_IFAR_WIDTH:61] cp_bp_t1_ifar,
   output [0:1]                cp_bp_t1_bh0_hist,
   output [0:1]                cp_bp_t1_bh1_hist,
   output [0:1]                cp_bp_t1_bh2_hist,
   output                      cp_bp_t1_br_pred,
   output                      cp_bp_t1_br_taken,
   output                      cp_bp_t1_bh_update,
   output                      cp_bp_t1_bcctr,
   output                      cp_bp_t1_bclr,
   output                      cp_bp_t1_getnia,
   output                      cp_bp_t1_group,
   output                      cp_bp_t1_lk,
   output [0:1]                cp_bp_t1_bh,
   output [0:9]                cp_bp_t1_gshare,
   output [0:2]                cp_bp_t1_ls_ptr,
   output [62-`EFF_IFAR_WIDTH:61] cp_bp_t1_ctr,
   output                      cp_bp_t1_btb_entry,
   output [0:1]                cp_bp_t1_btb_hist,
`endif

   // Output to dispatch to block due to ivax
   output [0:`THREADS-1]       cp_dis_ivax,

   // LQ Instruction Executed
   input [0:`THREADS-1]        lq0_iu_execute_vld,
   input [0:`ITAG_SIZE_ENC-1]  lq0_iu_itag,
   input                       lq0_iu_n_flush,
   input                       lq0_iu_np1_flush,
   input                       lq0_iu_dacr_type,
   input [0:3]                 lq0_iu_dacrw,
   input [0:31]                lq0_iu_instr,
   input [64-`GPR_WIDTH:63]    lq0_iu_eff_addr,
   input                       lq0_iu_exception_val,
   input [0:5]                 lq0_iu_exception,
   input                       lq0_iu_flush2ucode,
   input                       lq0_iu_flush2ucode_type,
   input [0:`THREADS-1]        lq0_iu_recirc_val,
   input [0:`THREADS-1]        lq0_iu_dear_val,

   input [0:`THREADS-1]        lq1_iu_execute_vld,
   input [0:`ITAG_SIZE_ENC-1]  lq1_iu_itag,
   input                       lq1_iu_n_flush,
   input                       lq1_iu_np1_flush,
   input                       lq1_iu_exception_val,
   input [0:5]                 lq1_iu_exception,
   input                       lq1_iu_dacr_type,
   input [0:3]                 lq1_iu_dacrw,
   input [0:3]                 lq1_iu_perf_events,

   output [0:`THREADS-1]       iu_lq_i0_completed,
   output [0:`THREADS-1]       iu_lq_i1_completed,
   output [0:`ITAG_SIZE_ENC-1] iu_lq_t0_i0_completed_itag,
   output [0:`ITAG_SIZE_ENC-1] iu_lq_t0_i1_completed_itag,
`ifndef THREADS1
   output [0:`ITAG_SIZE_ENC-1] iu_lq_t1_i0_completed_itag,
   output [0:`ITAG_SIZE_ENC-1] iu_lq_t1_i1_completed_itag,
`endif

   output [0:`THREADS-1]       iu_lq_recirc_val,

   // BR Instruction Executed
   input [0:`THREADS-1]        br_iu_execute_vld,
   input [0:`ITAG_SIZE_ENC-1]  br_iu_itag,
   input [0:`THREADS-1]        br_iu_redirect,
   input [62-`EFF_IFAR_ARCH:61] br_iu_bta,
   input                       br_iu_taken,
   input [0:3]                 br_iu_perf_events,

   // XU0 Instruction Executed
   input [0:`THREADS-1]        xu_iu_execute_vld,
   input [0:`ITAG_SIZE_ENC-1]  xu_iu_itag,
   input                       xu_iu_n_flush,
   input                       xu_iu_np1_flush,
   input                       xu_iu_flush2ucode,
   input                       xu_iu_exception_val,
   input [0:4]                 xu_iu_exception,
   input [0:`THREADS-1]        xu_iu_mtiar,
   input [62-`EFF_IFAR_ARCH:61] xu_iu_bta,
   input [0:3]                 xu_iu_perf_events,

   // XU0 Instruction Executed
   input [0:`THREADS-1]        xu1_iu_execute_vld,
   input [0:`ITAG_SIZE_ENC-1]  xu1_iu_itag,

   // AXU0 Instruction Executed
   input [0:`THREADS-1]        axu0_iu_execute_vld,
   input [0:`ITAG_SIZE_ENC-1]  axu0_iu_itag,
   input                       axu0_iu_n_flush,
   input                       axu0_iu_np1_flush,
   input                       axu0_iu_n_np1_flush,
   input                       axu0_iu_flush2ucode,
   input                       axu0_iu_flush2ucode_type,
   input                       axu0_iu_exception_val,
   input [0:3]                 axu0_iu_exception,
   input [0:3]                 axu0_iu_perf_events,

   // AXU1 Instruction Executed
   input [0:`THREADS-1]        axu1_iu_execute_vld,
   input [0:`ITAG_SIZE_ENC-1]  axu1_iu_itag,
   input                       axu1_iu_n_flush,
   input                       axu1_iu_np1_flush,
   input                       axu1_iu_flush2ucode,
   input                       axu1_iu_flush2ucode_type,
   input                       axu1_iu_exception_val,
   input [0:3]                 axu1_iu_exception,
   input [0:3]                 axu1_iu_perf_events,

   // Interrupts
	input [0:`THREADS-1]        an_ac_uncond_dbg_event,
   input [0:`THREADS-1]        xu_iu_external_mchk,
   input [0:`THREADS-1]        xu_iu_ext_interrupt,
   input [0:`THREADS-1]        xu_iu_dec_interrupt,
   input [0:`THREADS-1]        xu_iu_udec_interrupt,
   input [0:`THREADS-1]        xu_iu_perf_interrupt,
   input [0:`THREADS-1]        xu_iu_fit_interrupt,
   input [0:`THREADS-1]        xu_iu_crit_interrupt,
   input [0:`THREADS-1]        xu_iu_wdog_interrupt,
   input [0:`THREADS-1]        xu_iu_gwdog_interrupt,
   input [0:`THREADS-1]        xu_iu_gfit_interrupt,
   input [0:`THREADS-1]        xu_iu_gdec_interrupt,
   input [0:`THREADS-1]        xu_iu_dbell_interrupt,
   input [0:`THREADS-1]        xu_iu_cdbell_interrupt,
   input [0:`THREADS-1]        xu_iu_gdbell_interrupt,
   input [0:`THREADS-1]        xu_iu_gcdbell_interrupt,
   input [0:`THREADS-1]        xu_iu_gmcdbell_interrupt,
   input [0:`THREADS-1]        xu_iu_dbsr_ide,
   input [62-`EFF_IFAR_ARCH:61] xu_iu_t0_rest_ifar,
`ifndef THREADS1
   input [62-`EFF_IFAR_ARCH:61] xu_iu_t1_rest_ifar,
`endif
   input [0:`THREADS-1]        axu0_iu_async_fex,

   // To Ierats
   output                      cp_is_isync,		// Or together from each completion unit
   output                      cp_is_csync,		// Or together from each completion unit

   // Flushes
   output [0:`THREADS-1]       iu_flush,
   output [0:`THREADS-1]       cp_flush_into_uc,
   output [43:61]              cp_uc_t0_flush_ifar,
`ifndef THREADS1
   output [43:61]              cp_uc_t1_flush_ifar,
`endif
   output [0:`THREADS-1]       cp_uc_np1_flush,
   output [0:`THREADS-1]       cp_flush,
   output [0:`ITAG_SIZE_ENC-1]   cp_t0_next_itag,
   output [0:`ITAG_SIZE_ENC-1]   cp_t0_flush_itag,
   output [62-`EFF_IFAR_ARCH:61] cp_t0_flush_ifar,
`ifndef THREADS1
   output [0:`ITAG_SIZE_ENC-1]   cp_t1_next_itag,
   output [0:`ITAG_SIZE_ENC-1]   cp_t1_flush_itag,
   output [62-`EFF_IFAR_ARCH:61] cp_t1_flush_ifar,
`endif
   output [0:`THREADS-1]       cp_iu0_flush_2ucode,
   output [0:`THREADS-1]       cp_iu0_flush_2ucode_type,
   output [0:`THREADS-1]       cp_iu0_flush_nonspec,
   input                       pc_iu_init_reset,
   output [0:`THREADS-1]       cp_rn_uc_credit_free,

   // Signals to SPR partition
   output [0:`THREADS-1]       iu_xu_rfi,
   output [0:`THREADS-1]       iu_xu_rfgi,
   output [0:`THREADS-1]       iu_xu_rfci,
   output [0:`THREADS-1]       iu_xu_rfmci,
   output [0:`THREADS-1]       iu_xu_int,
   output [0:`THREADS-1]       iu_xu_gint,
   output [0:`THREADS-1]       iu_xu_cint,
   output [0:`THREADS-1]       iu_xu_mcint,
   output [0:`THREADS-1]       iu_xu_dear_update,
   output [0:`THREADS-1]       iu_spr_eheir_update,
   output [62-`EFF_IFAR_ARCH:61] iu_xu_t0_nia,
   output [0:16]               iu_xu_t0_esr,
   output [0:14]               iu_xu_t0_mcsr,
   output [0:18]               iu_xu_t0_dbsr,
   output [64-`GPR_WIDTH:63]   iu_xu_t0_dear,
   output [0:31]               iu_spr_t0_eheir,
   input [0:1]                 xu_iu_t0_dbcr0_dac1,
   input [0:1]                 xu_iu_t0_dbcr0_dac2,
   input [0:1]                 xu_iu_t0_dbcr0_dac3,
   input [0:1]                 xu_iu_t0_dbcr0_dac4,
`ifndef THREADS1
   output [62-`EFF_IFAR_ARCH:61] iu_xu_t1_nia,
   output [0:16]               iu_xu_t1_esr,
   output [0:14]               iu_xu_t1_mcsr,
   output [0:18]               iu_xu_t1_dbsr,
   output [64-`GPR_WIDTH:63]   iu_xu_t1_dear,
   output [0:31]               iu_spr_t1_eheir,
   input [0:1]                 xu_iu_t1_dbcr0_dac1,
   input [0:1]                 xu_iu_t1_dbcr0_dac2,
   input [0:1]                 xu_iu_t1_dbcr0_dac3,
   input [0:1]                 xu_iu_t1_dbcr0_dac4,
`endif
   output [0:`THREADS-1]       iu_xu_dbsr_update,
   output [0:`THREADS-1]       iu_xu_dbsr_ude,
   output [0:`THREADS-1]       iu_xu_dbsr_ide,
   output [0:`THREADS-1]       iu_xu_esr_update,
   output [0:`THREADS-1]       iu_xu_act,
   output [0:`THREADS-1]       iu_xu_dbell_taken,
   output [0:`THREADS-1]       iu_xu_cdbell_taken,
   output [0:`THREADS-1]       iu_xu_gdbell_taken,
   output [0:`THREADS-1]       iu_xu_gcdbell_taken,
   output [0:`THREADS-1]       iu_xu_gmcdbell_taken,
   output [0:`THREADS-1]       iu_xu_instr_cpl,
   input [0:`THREADS-1]        xu_iu_np1_async_flush,
   output [0:`THREADS-1]       iu_xu_async_complete,
   input [0:`THREADS-1]        dp_cp_hold_req,
   output [0:`THREADS-1]       iu_mm_hold_ack,
   input [0:`THREADS-1]        dp_cp_bus_snoop_hold_req,
   output [0:`THREADS-1]       iu_mm_bus_snoop_hold_ack,
   input [0:`THREADS-1]        xu_iu_msr_de,
   input [0:`THREADS-1]        xu_iu_msr_pr,
   input [0:`THREADS-1]        xu_iu_msr_cm,
   input [0:`THREADS-1]        xu_iu_msr_gs,
   input [0:`THREADS-1]        xu_iu_msr_me,
   input [0:`THREADS-1]        xu_iu_dbcr0_edm,
   input [0:`THREADS-1]        xu_iu_dbcr0_idm,
   input [0:`THREADS-1]        xu_iu_dbcr0_icmp,
   input [0:`THREADS-1]        xu_iu_dbcr0_brt,
   input [0:`THREADS-1]        xu_iu_dbcr0_irpt,
   input [0:`THREADS-1]        xu_iu_dbcr0_trap,
   input [0:`THREADS-1]        xu_iu_iac1_en,
   input [0:`THREADS-1]        xu_iu_iac2_en,
   input [0:`THREADS-1]        xu_iu_iac3_en,
   input [0:`THREADS-1]        xu_iu_iac4_en,
   input [0:`THREADS-1]        xu_iu_dbcr0_ret,
   input [0:`THREADS-1]        xu_iu_dbcr1_iac12m,
   input [0:`THREADS-1]        xu_iu_dbcr1_iac34m,
   input [0:`THREADS-1]        lq_iu_spr_dbcr3_ivc,
   input [0:`THREADS-1]        xu_iu_epcr_extgs,
   input [0:`THREADS-1]        xu_iu_epcr_dtlbgs,
   input [0:`THREADS-1]        xu_iu_epcr_itlbgs,
   input [0:`THREADS-1]        xu_iu_epcr_dsigs,
   input [0:`THREADS-1]        xu_iu_epcr_isigs,
   input [0:`THREADS-1]        xu_iu_epcr_duvd,
   input [0:`THREADS-1]        xu_iu_epcr_icm,
   input [0:`THREADS-1]        xu_iu_epcr_gicm,
   input                       xu_iu_spr_ccr2_en_dcr,
   input                       xu_iu_spr_ccr2_ucode_dis,
   input                       xu_iu_hid_mmu_mode,
   input                       xu_iu_xucr4_mmu_mchk,
   output [0:`THREADS-1]       iu_xu_quiesce,
   output [0:`THREADS-1]       iu_pc_quiesce,

   // MMU Errors
   input [0:`THREADS-1]        mm_iu_ierat_rel_val,
   input [0:`THREADS-1]        mm_iu_ierat_pt_fault,
   input [0:`THREADS-1]        mm_iu_ierat_lrat_miss,
   input [0:`THREADS-1]        mm_iu_ierat_tlb_inelig,
   input [0:`THREADS-1]        mm_iu_tlb_multihit_err,
   input [0:`THREADS-1]        mm_iu_tlb_par_err,
   input [0:`THREADS-1]        mm_iu_lru_par_err,
   input [0:`THREADS-1]        mm_iu_tlb_miss,
   input [0:`THREADS-1]        mm_iu_reload_hit,
   input [3:4]                 mm_iu_ierat_mmucr1,
   input [0:`THREADS-1]        ic_cp_nonspec_hit,


   output [0:5]                cp_mm_except_taken_t0,
`ifndef THREADS1
   output [0:5]                cp_mm_except_taken_t1,
`endif

   // SPRs
   input [0:`THREADS-1]        xu_iu_single_instr_mode,
   input [0:`THREADS-1]        spr_single_issue,
   input [64-`GPR_WIDTH:51]    spr_ivpr,
   input [64-`GPR_WIDTH:51]    spr_givpr,
   input [62-`EFF_IFAR_ARCH:61] spr_iac1,
   input [62-`EFF_IFAR_ARCH:61] spr_iac2,
   input [62-`EFF_IFAR_ARCH:61] spr_iac3,
   input [62-`EFF_IFAR_ARCH:61] spr_iac4,

   // XER read bus to RF for store conditionals
   output [0:`XER_POOL_ENC-1]  iu_rf_t0_xer_p,
`ifndef THREADS1
   output [0:`XER_POOL_ENC-1]  iu_rf_t1_xer_p,
`endif

   // Signals from pervasive
   input [0:`THREADS-1]        pc_iu_ram_active,
   input [0:`THREADS-1]        pc_iu_ram_flush_thread,
   input [0:`THREADS-1]        xu_iu_msrovride_enab,
   output                      iu_pc_ram_done,				// Need to Or these togther to create
   output                      iu_pc_ram_interrupt,		// Need to Or these togther to create
   output                      iu_pc_ram_unsupported,
   input [0:`THREADS-1]        pc_iu_stop,
   input [0:`THREADS-1]        pc_iu_step,
   input [0:2]                 pc_iu_t0_dbg_action,
`ifndef THREADS1
   input [0:2]                 pc_iu_t1_dbg_action,
`endif
   output [0:`THREADS-1]       iu_pc_step_done,
   output [0:`THREADS-1]       iu_pc_stop_dbg_event,
   output [0:`THREADS-1]       iu_pc_err_debug_event,
   output [0:`THREADS-1]       iu_pc_attention_instr,
   output [0:`THREADS-1]       iu_pc_err_mchk_disabled,
   output [0:`THREADS-1]       ac_an_debug_trigger,
   output [0:`THREADS-1]       iu_xu_stop,

   input                            pc_iu_trace_bus_enable,
   input [0:10]                     pc_iu_debug_mux_ctrls,
   input  [0:31]                    debug_bus_in,
   output [0:31]                    debug_bus_out,
   input  [0:3]                     coretrace_ctrls_in,
   output [0:3]                     coretrace_ctrls_out,


   // Power
   inout                       vdd,
   inout                       gnd);

   wire [0:`THREADS-1]          cp_is_isync_int;
   wire [0:`THREADS-1]          cp_is_csync_int;
   wire [0:`THREADS-1]          iu_pc_ram_done_int;
   wire [0:`THREADS-1]          iu_pc_ram_interrupt_int;
   wire [0:`THREADS-1]          iu_pc_ram_unsupported_int;

   wire [0:`THREADS-1]          iu_pc_stop_dbg_event_int[0:`THREADS-1];

   wire [0:31]                     unit_dbg_data0;
   wire [0:31]                     unit_dbg_data1;
   wire [0:31]                     unit_dbg_data2;
   wire [0:31]                     unit_dbg_data3;
   wire [0:31]                     unit_dbg_data4;
   wire [0:31]                     unit_dbg_data5;
   wire [0:31]                     unit_dbg_data6;
   wire [0:31]                     unit_dbg_data7;
   wire [0:31]                     unit_dbg_data8;
   wire [0:31]                     unit_dbg_data9;
   wire [0:31]                     unit_dbg_data10;
   wire [0:31]                     unit_dbg_data11;
   wire [0:31]                     unit_dbg_data12;
   wire [0:31]                     unit_dbg_data13;
   wire [0:31]                     unit_dbg_data14;
   wire [0:31]                     unit_dbg_data15;

   // for now assigning the debug to 0
   assign unit_dbg_data0  = 32'h00000000;
   assign unit_dbg_data1  = 32'h00000000;
   assign unit_dbg_data2  = 32'h00000000;
   assign unit_dbg_data3  = 32'h00000000;
   assign unit_dbg_data4  = 32'h00000000;
   assign unit_dbg_data5  = 32'h00000000;
   assign unit_dbg_data6  = 32'h00000000;
   assign unit_dbg_data7  = 32'h00000000;
   assign unit_dbg_data8  = 32'h00000000;
   assign unit_dbg_data9  = 32'h00000000;
   assign unit_dbg_data10 = 32'h00000000;
   assign unit_dbg_data11 = 32'h00000000;
   assign unit_dbg_data12 = 32'h00000000;
   assign unit_dbg_data13 = 32'h00000000;
   assign unit_dbg_data14 = 32'h00000000;
   assign unit_dbg_data15 = 32'h00000000;



   assign cp_is_isync = |cp_is_isync_int;
   assign cp_is_csync = |cp_is_csync_int;
   assign iu_pc_ram_done = |iu_pc_ram_done_int;
   assign iu_pc_ram_interrupt = |iu_pc_ram_interrupt_int;
   assign iu_pc_ram_unsupported = |iu_pc_ram_unsupported_int;
 `ifdef THREADS1
   assign iu_pc_stop_dbg_event = iu_pc_stop_dbg_event_int[0][0];
 `endif
 `ifndef THREADS1
   assign iu_pc_stop_dbg_event = {(iu_pc_stop_dbg_event_int[0][0] | iu_pc_stop_dbg_event_int[1][1]), (iu_pc_stop_dbg_event_int[0][1] | iu_pc_stop_dbg_event_int[1][0])};
 `endif

	iuq_cpl iuq_cpl0(
      .vdd(vdd),
      .gnd(gnd),
      .nclk(nclk),
      .tc_ac_ccflush_dc(tc_ac_ccflush_dc),
      .clkoff_dc_b(clkoff_dc_b),
      .d_mode_dc(d_mode_dc),
      .delay_lclkr_dc(delay_lclkr_dc),
      .mpw1_dc_b(mpw1_dc_b),
      .mpw2_dc_b(mpw2_dc_b),
      .func_sl_thold_2(pc_iu_func_sl_thold_2),
      .func_slp_sl_thold_2(pc_iu_func_slp_sl_thold_2),
      .sg_2(pc_iu_sg_2),
      .scan_in(cp_scan_in[0]),
      .scan_out(cp_scan_out[0]),
      .pc_iu_event_bus_enable(pc_iu_event_bus_enable),
      .pc_iu_event_count_mode(pc_iu_event_count_mode),
      .spr_cp_perf_event_mux_ctrls(spr_cp_perf_event_mux_ctrls[0:15]),
      .event_bus_in(event_bus_in[0:3]),
      .event_bus_out(event_bus_out[0:3]),
      .rn_cp_iu6_i0_vld(rn_cp_iu6_t0_i0_vld),
      .rn_cp_iu6_i0_itag(rn_cp_iu6_t0_i0_itag),
      .rn_cp_iu6_i0_ucode(rn_cp_iu6_t0_i0_ucode),
      .rn_cp_iu6_i0_fuse_nop(rn_cp_iu6_t0_i0_fuse_nop),
      .rn_cp_iu6_i0_rte_lq(rn_cp_iu6_t0_i0_rte_lq),
      .rn_cp_iu6_i0_rte_sq(rn_cp_iu6_t0_i0_rte_sq),
      .rn_cp_iu6_i0_rte_fx0(rn_cp_iu6_t0_i0_rte_fx0),
      .rn_cp_iu6_i0_rte_fx1(rn_cp_iu6_t0_i0_rte_fx1),
      .rn_cp_iu6_i0_rte_axu0(rn_cp_iu6_t0_i0_rte_axu0),
      .rn_cp_iu6_i0_rte_axu1(rn_cp_iu6_t0_i0_rte_axu1),
      .rn_cp_iu6_i0_ifar(rn_cp_iu6_t0_i0_ifar),
      .rn_cp_iu6_i0_bta(rn_cp_iu6_t0_i0_bta),
      .rn_cp_iu6_i0_isram(rn_cp_iu6_t0_i0_isram),
      .rn_cp_iu6_i0_instr(rn_cp_iu6_t0_i0_instr),
      .rn_cp_iu6_i0_valop(rn_cp_iu6_t0_i0_valop),
      .rn_cp_iu6_i0_error(rn_cp_iu6_t0_i0_error),
      .rn_cp_iu6_i0_br_pred(rn_cp_iu6_t0_i0_br_pred),
      .rn_cp_iu6_i0_bh_update(rn_cp_iu6_t0_i0_bh_update),
      .rn_cp_iu6_i0_bh0_hist(rn_cp_iu6_t0_i0_bh0_hist),
      .rn_cp_iu6_i0_bh1_hist(rn_cp_iu6_t0_i0_bh1_hist),
      .rn_cp_iu6_i0_bh2_hist(rn_cp_iu6_t0_i0_bh2_hist),
      .rn_cp_iu6_i0_gshare(rn_cp_iu6_t0_i0_gshare),
      .rn_cp_iu6_i0_ls_ptr(rn_cp_iu6_t0_i0_ls_ptr),
      .rn_cp_iu6_i0_match(rn_cp_iu6_t0_i0_match),
      .rn_cp_iu6_i0_type_fp(rn_cp_iu6_t0_i0_type_fp),
      .rn_cp_iu6_i0_type_ap(rn_cp_iu6_t0_i0_type_ap),
      .rn_cp_iu6_i0_type_spv(rn_cp_iu6_t0_i0_type_spv),
      .rn_cp_iu6_i0_type_st(rn_cp_iu6_t0_i0_type_st),
      .rn_cp_iu6_i0_async_block(rn_cp_iu6_t0_i0_async_block),
      .rn_cp_iu6_i0_np1_flush(rn_cp_iu6_t0_i0_np1_flush),
      .rn_cp_iu6_i0_t1_v(rn_cp_iu6_t0_i0_t1_v),
      .rn_cp_iu6_i0_t1_t(rn_cp_iu6_t0_i0_t1_t),
      .rn_cp_iu6_i0_t1_p(rn_cp_iu6_t0_i0_t1_p),
      .rn_cp_iu6_i0_t1_a(rn_cp_iu6_t0_i0_t1_a),
      .rn_cp_iu6_i0_t2_v(rn_cp_iu6_t0_i0_t2_v),
      .rn_cp_iu6_i0_t2_t(rn_cp_iu6_t0_i0_t2_t),
      .rn_cp_iu6_i0_t2_p(rn_cp_iu6_t0_i0_t2_p),
      .rn_cp_iu6_i0_t2_a(rn_cp_iu6_t0_i0_t2_a),
      .rn_cp_iu6_i0_t3_v(rn_cp_iu6_t0_i0_t3_v),
      .rn_cp_iu6_i0_t3_t(rn_cp_iu6_t0_i0_t3_t),
      .rn_cp_iu6_i0_t3_p(rn_cp_iu6_t0_i0_t3_p),
      .rn_cp_iu6_i0_t3_a(rn_cp_iu6_t0_i0_t3_a),
      .rn_cp_iu6_i0_btb_entry(rn_cp_iu6_t0_i0_btb_entry),
      .rn_cp_iu6_i0_btb_hist(rn_cp_iu6_t0_i0_btb_hist),
      .rn_cp_iu6_i0_bta_val(rn_cp_iu6_t0_i0_bta_val),
      .rn_cp_iu6_i1_vld(rn_cp_iu6_t0_i1_vld),
      .rn_cp_iu6_i1_itag(rn_cp_iu6_t0_i1_itag),
      .rn_cp_iu6_i1_ucode(rn_cp_iu6_t0_i1_ucode),
      .rn_cp_iu6_i1_fuse_nop(rn_cp_iu6_t0_i1_fuse_nop),
      .rn_cp_iu6_i1_rte_lq(rn_cp_iu6_t0_i1_rte_lq),
      .rn_cp_iu6_i1_rte_sq(rn_cp_iu6_t0_i1_rte_sq),
      .rn_cp_iu6_i1_rte_fx0(rn_cp_iu6_t0_i1_rte_fx0),
      .rn_cp_iu6_i1_rte_fx1(rn_cp_iu6_t0_i1_rte_fx1),
      .rn_cp_iu6_i1_rte_axu0(rn_cp_iu6_t0_i1_rte_axu0),
      .rn_cp_iu6_i1_rte_axu1(rn_cp_iu6_t0_i1_rte_axu1),
      .rn_cp_iu6_i1_ifar(rn_cp_iu6_t0_i1_ifar),
      .rn_cp_iu6_i1_bta(rn_cp_iu6_t0_i1_bta),
      .rn_cp_iu6_i1_isram(rn_cp_iu6_t0_i1_isram),
      .rn_cp_iu6_i1_instr(rn_cp_iu6_t0_i1_instr),
      .rn_cp_iu6_i1_valop(rn_cp_iu6_t0_i1_valop),
      .rn_cp_iu6_i1_error(rn_cp_iu6_t0_i1_error),
      .rn_cp_iu6_i1_br_pred(rn_cp_iu6_t0_i1_br_pred),
      .rn_cp_iu6_i1_bh_update(rn_cp_iu6_t0_i1_bh_update),
      .rn_cp_iu6_i1_bh0_hist(rn_cp_iu6_t0_i1_bh0_hist),
      .rn_cp_iu6_i1_bh1_hist(rn_cp_iu6_t0_i1_bh1_hist),
      .rn_cp_iu6_i1_bh2_hist(rn_cp_iu6_t0_i1_bh2_hist),
      .rn_cp_iu6_i1_gshare(rn_cp_iu6_t0_i1_gshare),
      .rn_cp_iu6_i1_ls_ptr(rn_cp_iu6_t0_i1_ls_ptr),
      .rn_cp_iu6_i1_match(rn_cp_iu6_t0_i1_match),
      .rn_cp_iu6_i1_type_fp(rn_cp_iu6_t0_i1_type_fp),
      .rn_cp_iu6_i1_type_ap(rn_cp_iu6_t0_i1_type_ap),
      .rn_cp_iu6_i1_type_spv(rn_cp_iu6_t0_i1_type_spv),
      .rn_cp_iu6_i1_type_st(rn_cp_iu6_t0_i1_type_st),
      .rn_cp_iu6_i1_async_block(rn_cp_iu6_t0_i1_async_block),
      .rn_cp_iu6_i1_np1_flush(rn_cp_iu6_t0_i1_np1_flush),
      .rn_cp_iu6_i1_t1_v(rn_cp_iu6_t0_i1_t1_v),
      .rn_cp_iu6_i1_t1_t(rn_cp_iu6_t0_i1_t1_t),
      .rn_cp_iu6_i1_t1_p(rn_cp_iu6_t0_i1_t1_p),
      .rn_cp_iu6_i1_t1_a(rn_cp_iu6_t0_i1_t1_a),
      .rn_cp_iu6_i1_t2_v(rn_cp_iu6_t0_i1_t2_v),
      .rn_cp_iu6_i1_t2_t(rn_cp_iu6_t0_i1_t2_t),
      .rn_cp_iu6_i1_t2_p(rn_cp_iu6_t0_i1_t2_p),
      .rn_cp_iu6_i1_t2_a(rn_cp_iu6_t0_i1_t2_a),
      .rn_cp_iu6_i1_t3_v(rn_cp_iu6_t0_i1_t3_v),
      .rn_cp_iu6_i1_t3_t(rn_cp_iu6_t0_i1_t3_t),
      .rn_cp_iu6_i1_t3_p(rn_cp_iu6_t0_i1_t3_p),
      .rn_cp_iu6_i1_t3_a(rn_cp_iu6_t0_i1_t3_a),
      .rn_cp_iu6_i1_btb_entry(rn_cp_iu6_t0_i1_btb_entry),
      .rn_cp_iu6_i1_btb_hist(rn_cp_iu6_t0_i1_btb_hist),
      .rn_cp_iu6_i1_bta_val(rn_cp_iu6_t0_i1_bta_val),
      .cp_rn_empty(cp_rn_empty[0]),
      .cp_async_block(cp_async_block[0]),
      .cp_rn_i0_v(cp_rn_t0_i0_v),
      .cp_rn_i0_axu_exception_val(cp_rn_t0_i0_axu_exception_val),
      .cp_rn_i0_axu_exception(cp_rn_t0_i0_axu_exception),
      .cp_rn_i0_t1_v(cp_rn_t0_i0_t1_v),
      .cp_rn_i0_t1_t(cp_rn_t0_i0_t1_t),
      .cp_rn_i0_t1_p(cp_rn_t0_i0_t1_p),
      .cp_rn_i0_t1_a(cp_rn_t0_i0_t1_a),
      .cp_rn_i0_t2_v(cp_rn_t0_i0_t2_v),
      .cp_rn_i0_t2_t(cp_rn_t0_i0_t2_t),
      .cp_rn_i0_t2_p(cp_rn_t0_i0_t2_p),
      .cp_rn_i0_t2_a(cp_rn_t0_i0_t2_a),
      .cp_rn_i0_t3_v(cp_rn_t0_i0_t3_v),
      .cp_rn_i0_t3_t(cp_rn_t0_i0_t3_t),
      .cp_rn_i0_t3_p(cp_rn_t0_i0_t3_p),
      .cp_rn_i0_t3_a(cp_rn_t0_i0_t3_a),
      .cp_rn_i1_v(cp_rn_t0_i1_v),
      .cp_rn_i1_axu_exception_val(cp_rn_t0_i1_axu_exception_val),
      .cp_rn_i1_axu_exception(cp_rn_t0_i1_axu_exception),
      .cp_rn_i1_t1_v(cp_rn_t0_i1_t1_v),
      .cp_rn_i1_t1_t(cp_rn_t0_i1_t1_t),
      .cp_rn_i1_t1_p(cp_rn_t0_i1_t1_p),
      .cp_rn_i1_t1_a(cp_rn_t0_i1_t1_a),
      .cp_rn_i1_t2_v(cp_rn_t0_i1_t2_v),
      .cp_rn_i1_t2_t(cp_rn_t0_i1_t2_t),
      .cp_rn_i1_t2_p(cp_rn_t0_i1_t2_p),
      .cp_rn_i1_t2_a(cp_rn_t0_i1_t2_a),
      .cp_rn_i1_t3_v(cp_rn_t0_i1_t3_v),
      .cp_rn_i1_t3_t(cp_rn_t0_i1_t3_t),
      .cp_rn_i1_t3_p(cp_rn_t0_i1_t3_p),
      .cp_rn_i1_t3_a(cp_rn_t0_i1_t3_a),
      .cp_bp_val(cp_bp_t0_val),
      .cp_bp_ifar(cp_bp_t0_ifar),
      .cp_bp_bh0_hist(cp_bp_t0_bh0_hist),
      .cp_bp_bh1_hist(cp_bp_t0_bh1_hist),
      .cp_bp_bh2_hist(cp_bp_t0_bh2_hist),
      .cp_bp_br_pred(cp_bp_t0_br_pred),
      .cp_bp_br_taken(cp_bp_t0_br_taken),
      .cp_bp_bh_update(cp_bp_t0_bh_update),
      .cp_bp_bcctr(cp_bp_t0_bcctr),
      .cp_bp_bclr(cp_bp_t0_bclr),
      .cp_bp_getnia(cp_bp_t0_getnia),
      .cp_bp_group(cp_bp_t0_group),
      .cp_dis_ivax(cp_dis_ivax[0]),
      .cp_bp_lk(cp_bp_t0_lk),
      .cp_bp_bh(cp_bp_t0_bh),
      .cp_bp_gshare(cp_bp_t0_gshare),
      .cp_bp_ls_ptr(cp_bp_t0_ls_ptr),
      .cp_bp_ctr(cp_bp_t0_ctr),
      .cp_bp_btb_entry(cp_bp_t0_btb_entry),
      .cp_bp_btb_hist(cp_bp_t0_btb_hist),
      .lq0_iu_execute_vld(lq0_iu_execute_vld[0]),
      .lq0_iu_itag(lq0_iu_itag),
      .lq0_iu_n_flush(lq0_iu_n_flush),
      .lq0_iu_np1_flush(lq0_iu_np1_flush),
      .lq0_iu_dacr_type(lq0_iu_dacr_type),
      .lq0_iu_dacrw(lq0_iu_dacrw),
      .lq0_iu_instr(lq0_iu_instr),
      .lq0_iu_eff_addr(lq0_iu_eff_addr),
      .lq0_iu_exception_val(lq0_iu_exception_val),
      .lq0_iu_exception(lq0_iu_exception),
      .lq0_iu_flush2ucode(lq0_iu_flush2ucode),
      .lq0_iu_flush2ucode_type(lq0_iu_flush2ucode_type),
      .lq0_iu_recirc_val(lq0_iu_recirc_val[0]),
      .lq0_iu_dear_val(lq0_iu_dear_val[0]),
      .lq1_iu_execute_vld(lq1_iu_execute_vld[0]),
      .lq1_iu_itag(lq1_iu_itag),
      .lq1_iu_n_flush(lq1_iu_n_flush),
      .lq1_iu_np1_flush(lq1_iu_np1_flush),
      .lq1_iu_exception_val(lq1_iu_exception_val),
      .lq1_iu_exception(lq1_iu_exception),
      .lq1_iu_dacr_type(lq1_iu_dacr_type),
      .lq1_iu_dacrw(lq1_iu_dacrw),
      .lq1_iu_perf_events(lq1_iu_perf_events),
      .iu_lq_i0_completed(iu_lq_i0_completed[0]),
      .iu_lq_i1_completed(iu_lq_i1_completed[0]),
      .iu_lq_i0_completed_itag(iu_lq_t0_i0_completed_itag),
      .iu_lq_i1_completed_itag(iu_lq_t0_i1_completed_itag),
      .iu_lq_recirc_val(iu_lq_recirc_val[0]),
      .br_iu_execute_vld(br_iu_execute_vld[0]),
      .br_iu_itag(br_iu_itag),
      .br_iu_bta(br_iu_bta),
      .br_iu_redirect(br_iu_redirect[0]),
      .br_iu_taken(br_iu_taken),
      .br_iu_perf_events(br_iu_perf_events),
      .xu_iu_execute_vld(xu_iu_execute_vld[0]),
      .xu_iu_itag(xu_iu_itag),
      .xu_iu_exception_val(xu_iu_exception_val),
      .xu_iu_exception(xu_iu_exception),
      .xu_iu_mtiar(xu_iu_mtiar[0]),
      .xu_iu_bta(xu_iu_bta),
      .xu_iu_perf_events(xu_iu_perf_events),
      .xu_iu_n_flush(xu_iu_n_flush),
      .xu_iu_np1_flush(xu_iu_np1_flush),
      .xu_iu_flush2ucode(xu_iu_flush2ucode),
      .xu1_iu_execute_vld(xu1_iu_execute_vld[0]),
      .xu1_iu_itag(xu1_iu_itag),
      .axu0_iu_execute_vld(axu0_iu_execute_vld[0]),
      .axu0_iu_itag(axu0_iu_itag),
      .axu0_iu_n_flush(axu0_iu_n_flush),
      .axu0_iu_np1_flush(axu0_iu_np1_flush),
      .axu0_iu_n_np1_flush(axu0_iu_n_np1_flush),
      .axu0_iu_exception(axu0_iu_exception),
      .axu0_iu_exception_val(axu0_iu_exception_val),
      .axu0_iu_flush2ucode(axu0_iu_flush2ucode),
      .axu0_iu_flush2ucode_type(axu0_iu_flush2ucode_type),
      .axu0_iu_async_fex(axu0_iu_async_fex[0]),
      .axu0_iu_perf_events(axu0_iu_perf_events),
      .axu1_iu_execute_vld(axu1_iu_execute_vld[0]),
      .axu1_iu_itag(axu1_iu_itag),
      .axu1_iu_n_flush(axu1_iu_n_flush),
      .axu1_iu_np1_flush(axu1_iu_np1_flush),
      .axu1_iu_exception(axu1_iu_exception),
      .axu1_iu_exception_val(axu1_iu_exception_val),
      .axu1_iu_flush2ucode(axu1_iu_flush2ucode),
      .axu1_iu_flush2ucode_type(axu1_iu_flush2ucode_type),
      .axu1_iu_perf_events(axu1_iu_perf_events),
      .an_ac_uncond_dbg_event(an_ac_uncond_dbg_event[0]),
      .xu_iu_external_mchk(xu_iu_external_mchk[0]),
      .xu_iu_ext_interrupt(xu_iu_ext_interrupt[0]),
      .xu_iu_dec_interrupt(xu_iu_dec_interrupt[0]),
      .xu_iu_udec_interrupt(xu_iu_udec_interrupt[0]),
      .xu_iu_perf_interrupt(xu_iu_perf_interrupt[0]),
      .xu_iu_fit_interrupt(xu_iu_fit_interrupt[0]),
      .xu_iu_crit_interrupt(xu_iu_crit_interrupt[0]),
      .xu_iu_wdog_interrupt(xu_iu_wdog_interrupt[0]),
      .xu_iu_gwdog_interrupt(xu_iu_gwdog_interrupt[0]),
      .xu_iu_gfit_interrupt(xu_iu_gfit_interrupt[0]),
      .xu_iu_gdec_interrupt(xu_iu_gdec_interrupt[0]),
      .xu_iu_dbell_interrupt(xu_iu_dbell_interrupt[0]),
      .xu_iu_cdbell_interrupt(xu_iu_cdbell_interrupt[0]),
      .xu_iu_gdbell_interrupt(xu_iu_gdbell_interrupt[0]),
      .xu_iu_gcdbell_interrupt(xu_iu_gcdbell_interrupt[0]),
      .xu_iu_gmcdbell_interrupt(xu_iu_gmcdbell_interrupt[0]),
      .xu_iu_dbsr_ide(xu_iu_dbsr_ide[0]),
      .xu_iu_rest_ifar(xu_iu_t0_rest_ifar),
      .cp_is_isync(cp_is_isync_int[0]),
      .cp_is_csync(cp_is_csync_int[0]),
      .iu_flush(iu_flush[0]),
      .cp_flush_into_uc(cp_flush_into_uc[0]),
      .cp_uc_flush_ifar(cp_uc_t0_flush_ifar),
      .cp_uc_np1_flush(cp_uc_np1_flush[0]),
      .cp_flush(cp_flush[0]),
      .cp_next_itag(cp_t0_next_itag),
      .cp_flush_itag(cp_t0_flush_itag),
      .cp_flush_ifar(cp_t0_flush_ifar),
      .cp_iu0_flush_2ucode(cp_iu0_flush_2ucode[0]),
      .cp_iu0_flush_2ucode_type(cp_iu0_flush_2ucode_type[0]),
      .cp_iu0_flush_nonspec(cp_iu0_flush_nonspec[0]),
      .pc_iu_init_reset(pc_iu_init_reset),
      .cp_rn_uc_credit_free(cp_rn_uc_credit_free[0]),
      .iu_xu_rfi(iu_xu_rfi[0]),
      .iu_xu_rfgi(iu_xu_rfgi[0]),
      .iu_xu_rfci(iu_xu_rfci[0]),
      .iu_xu_rfmci(iu_xu_rfmci[0]),
      .iu_xu_int(iu_xu_int[0]),
      .iu_xu_gint(iu_xu_gint[0]),
      .iu_xu_cint(iu_xu_cint[0]),
      .iu_xu_mcint(iu_xu_mcint[0]),
      .iu_xu_nia(iu_xu_t0_nia),
      .iu_xu_esr(iu_xu_t0_esr),
      .iu_xu_mcsr(iu_xu_t0_mcsr),
      .iu_xu_dbsr(iu_xu_t0_dbsr),
      .iu_xu_dear_update(iu_xu_dear_update[0]),
      .iu_xu_dear(iu_xu_t0_dear),
      .iu_xu_dbsr_update(iu_xu_dbsr_update[0]),
      .iu_xu_dbsr_ude(iu_xu_dbsr_ude[0]),
      .iu_xu_dbsr_ide(iu_xu_dbsr_ide[0]),
      .iu_xu_esr_update(iu_xu_esr_update[0]),
      .iu_xu_act(iu_xu_act[0]),
      .iu_xu_dbell_taken(iu_xu_dbell_taken[0]),
      .iu_xu_cdbell_taken(iu_xu_cdbell_taken[0]),
      .iu_xu_gdbell_taken(iu_xu_gdbell_taken[0]),
      .iu_xu_gcdbell_taken(iu_xu_gcdbell_taken[0]),
      .iu_xu_gmcdbell_taken(iu_xu_gmcdbell_taken[0]),
      .iu_xu_instr_cpl(iu_xu_instr_cpl[0]),
      .xu_iu_np1_async_flush(xu_iu_np1_async_flush[0]),
      .iu_xu_async_complete(iu_xu_async_complete[0]),
      .dp_cp_hold_req(dp_cp_hold_req[0]),
      .iu_mm_hold_ack(iu_mm_hold_ack[0]),
      .dp_cp_bus_snoop_hold_req(dp_cp_bus_snoop_hold_req[0]),
      .iu_mm_bus_snoop_hold_ack(iu_mm_bus_snoop_hold_ack[0]),
      .iu_spr_eheir_update(iu_spr_eheir_update[0]),
      .iu_spr_eheir(iu_spr_t0_eheir),
      .xu_iu_msr_de(xu_iu_msr_de[0]),
      .xu_iu_msr_pr(xu_iu_msr_pr[0]),
      .xu_iu_msr_cm(xu_iu_msr_cm[0]),
      .xu_iu_msr_gs(xu_iu_msr_gs[0]),
      .xu_iu_msr_me(xu_iu_msr_me[0]),
      .xu_iu_dbcr0_edm(xu_iu_dbcr0_edm[0]),
      .xu_iu_dbcr0_idm(xu_iu_dbcr0_idm[0]),
      .xu_iu_dbcr0_icmp(xu_iu_dbcr0_icmp[0]),
      .xu_iu_dbcr0_brt(xu_iu_dbcr0_brt[0]),
      .xu_iu_dbcr0_irpt(xu_iu_dbcr0_irpt[0]),
      .xu_iu_dbcr0_trap(xu_iu_dbcr0_trap[0]),
      .xu_iu_iac1_en(xu_iu_iac1_en[0]),
      .xu_iu_iac2_en(xu_iu_iac2_en[0]),
      .xu_iu_iac3_en(xu_iu_iac3_en[0]),
      .xu_iu_iac4_en(xu_iu_iac4_en[0]),
      .xu_iu_dbcr0_dac1(xu_iu_t0_dbcr0_dac1),
      .xu_iu_dbcr0_dac2(xu_iu_t0_dbcr0_dac2),
      .xu_iu_dbcr0_dac3(xu_iu_t0_dbcr0_dac3),
      .xu_iu_dbcr0_dac4(xu_iu_t0_dbcr0_dac4),
      .xu_iu_dbcr0_ret(xu_iu_dbcr0_ret[0]),
      .xu_iu_dbcr1_iac12m(xu_iu_dbcr1_iac12m[0]),
      .xu_iu_dbcr1_iac34m(xu_iu_dbcr1_iac34m[0]),
      .lq_iu_spr_dbcr3_ivc(lq_iu_spr_dbcr3_ivc[0]),
      .xu_iu_epcr_extgs(xu_iu_epcr_extgs[0]),
      .xu_iu_epcr_dtlbgs(xu_iu_epcr_dtlbgs[0]),
      .xu_iu_epcr_itlbgs(xu_iu_epcr_itlbgs[0]),
      .xu_iu_epcr_dsigs(xu_iu_epcr_dsigs[0]),
      .xu_iu_epcr_isigs(xu_iu_epcr_isigs[0]),
      .xu_iu_epcr_duvd(xu_iu_epcr_duvd[0]),
      .xu_iu_epcr_icm(xu_iu_epcr_icm[0]),
      .xu_iu_epcr_gicm(xu_iu_epcr_gicm[0]),
      .xu_iu_ccr2_en_dcr(xu_iu_spr_ccr2_en_dcr),
      .xu_iu_ccr2_ucode_dis(xu_iu_spr_ccr2_ucode_dis),
      .xu_iu_hid_mmu_mode(xu_iu_hid_mmu_mode),
      .xu_iu_xucr4_mmu_mchk(xu_iu_xucr4_mmu_mchk),
      .iu_xu_quiesce(iu_xu_quiesce[0]),
      .iu_pc_quiesce(iu_pc_quiesce[0]),
      .mm_iu_ierat_rel_val(mm_iu_ierat_rel_val[0]),
      .mm_iu_ierat_pt_fault(mm_iu_ierat_pt_fault[0]),
      .mm_iu_ierat_lrat_miss(mm_iu_ierat_lrat_miss[0]),
      .mm_iu_ierat_tlb_inelig(mm_iu_ierat_tlb_inelig[0]),
      .mm_iu_tlb_multihit_err(mm_iu_tlb_multihit_err[0]),
      .mm_iu_tlb_par_err(mm_iu_tlb_par_err[0]),
      .mm_iu_lru_par_err(mm_iu_lru_par_err[0]),
      .mm_iu_tlb_miss(mm_iu_tlb_miss[0]),
      .mm_iu_reload_hit(mm_iu_reload_hit[0]),
      .mm_iu_ierat_mmucr1(mm_iu_ierat_mmucr1[3:4]),
      .ic_cp_nonspec_hit(ic_cp_nonspec_hit[0]),
      .cp_mm_except_taken(cp_mm_except_taken_t0),
      .xu_iu_single_instr_mode(xu_iu_single_instr_mode[0]),
      .spr_single_issue(spr_single_issue[0]),
      .spr_ivpr(spr_ivpr),
      .spr_givpr(spr_givpr),
      .spr_iac1(spr_iac1),
      .spr_iac2(spr_iac2),
      .spr_iac3(spr_iac3),
      .spr_iac4(spr_iac4),
      .iu_rf_xer_p(iu_rf_t0_xer_p),
      .pc_iu_ram_active(pc_iu_ram_active[0]),
      .pc_iu_ram_flush_thread(pc_iu_ram_flush_thread[0]),
      .xu_iu_msrovride_enab(xu_iu_msrovride_enab[0]),
      .iu_pc_ram_done(iu_pc_ram_done_int[0]),
      .iu_pc_ram_interrupt(iu_pc_ram_interrupt_int[0]),
      .iu_pc_ram_unsupported(iu_pc_ram_unsupported_int[0]),
      .pc_iu_stop(pc_iu_stop[0]),
      .pc_iu_step(pc_iu_step[0]),
      .pc_iu_dbg_action(pc_iu_t0_dbg_action),
      .iu_pc_step_done(iu_pc_step_done[0]),
      .iu_pc_stop_dbg_event(iu_pc_stop_dbg_event_int[0]),
      .iu_pc_err_debug_event(iu_pc_err_debug_event[0]),
      .iu_pc_attention_instr(iu_pc_attention_instr[0]),
      .iu_pc_err_mchk_disabled(iu_pc_err_mchk_disabled[0]),
      .ac_an_debug_trigger(ac_an_debug_trigger[0]),
      .iu_xu_stop(iu_xu_stop[0])
   );

`ifndef THREADS1
	iuq_cpl iuq_cpl1(
      .vdd(vdd),
      .gnd(gnd),
      .nclk(nclk),
      .tc_ac_ccflush_dc(tc_ac_ccflush_dc),
      .clkoff_dc_b(clkoff_dc_b),
      .d_mode_dc(d_mode_dc),
      .delay_lclkr_dc(delay_lclkr_dc),
      .mpw1_dc_b(mpw1_dc_b),
      .mpw2_dc_b(mpw2_dc_b),
      .func_sl_thold_2(pc_iu_func_sl_thold_2),
      .func_slp_sl_thold_2(pc_iu_func_slp_sl_thold_2),
      .sg_2(pc_iu_sg_2),
      .scan_in(cp_scan_in[1]),
      .scan_out(cp_scan_out[1]),
      .pc_iu_event_bus_enable(pc_iu_event_bus_enable),
      .pc_iu_event_count_mode(pc_iu_event_count_mode),
      .spr_cp_perf_event_mux_ctrls(spr_cp_perf_event_mux_ctrls[16:31]),
      .event_bus_in(event_bus_in[4:7]),
      .event_bus_out(event_bus_out[4:7]),
      .rn_cp_iu6_i0_vld(rn_cp_iu6_t1_i0_vld),
      .rn_cp_iu6_i0_itag(rn_cp_iu6_t1_i0_itag),
      .rn_cp_iu6_i0_ucode(rn_cp_iu6_t1_i0_ucode),
      .rn_cp_iu6_i0_fuse_nop(rn_cp_iu6_t1_i0_fuse_nop),
      .rn_cp_iu6_i0_rte_lq(rn_cp_iu6_t1_i0_rte_lq),
      .rn_cp_iu6_i0_rte_sq(rn_cp_iu6_t1_i0_rte_sq),
      .rn_cp_iu6_i0_rte_fx0(rn_cp_iu6_t1_i0_rte_fx0),
      .rn_cp_iu6_i0_rte_fx1(rn_cp_iu6_t1_i0_rte_fx1),
      .rn_cp_iu6_i0_rte_axu0(rn_cp_iu6_t1_i0_rte_axu0),
      .rn_cp_iu6_i0_rte_axu1(rn_cp_iu6_t1_i0_rte_axu1),
      .rn_cp_iu6_i0_ifar(rn_cp_iu6_t1_i0_ifar),
      .rn_cp_iu6_i0_bta(rn_cp_iu6_t1_i0_bta),
      .rn_cp_iu6_i0_isram(rn_cp_iu6_t1_i0_isram),
      .rn_cp_iu6_i0_instr(rn_cp_iu6_t1_i0_instr),
      .rn_cp_iu6_i0_valop(rn_cp_iu6_t1_i0_valop),
      .rn_cp_iu6_i0_error(rn_cp_iu6_t1_i0_error),
      .rn_cp_iu6_i0_br_pred(rn_cp_iu6_t1_i0_br_pred),
      .rn_cp_iu6_i0_bh_update(rn_cp_iu6_t1_i0_bh_update),
      .rn_cp_iu6_i0_bh0_hist(rn_cp_iu6_t1_i0_bh0_hist),
      .rn_cp_iu6_i0_bh1_hist(rn_cp_iu6_t1_i0_bh1_hist),
      .rn_cp_iu6_i0_bh2_hist(rn_cp_iu6_t1_i0_bh2_hist),
      .rn_cp_iu6_i0_gshare(rn_cp_iu6_t1_i0_gshare),
      .rn_cp_iu6_i0_ls_ptr(rn_cp_iu6_t1_i0_ls_ptr),
      .rn_cp_iu6_i0_match(rn_cp_iu6_t1_i0_match),
      .rn_cp_iu6_i0_type_fp(rn_cp_iu6_t1_i0_type_fp),
      .rn_cp_iu6_i0_type_ap(rn_cp_iu6_t1_i0_type_ap),
      .rn_cp_iu6_i0_type_spv(rn_cp_iu6_t1_i0_type_spv),
      .rn_cp_iu6_i0_type_st(rn_cp_iu6_t1_i0_type_st),
      .rn_cp_iu6_i0_async_block(rn_cp_iu6_t1_i0_async_block),
      .rn_cp_iu6_i0_np1_flush(rn_cp_iu6_t1_i0_np1_flush),
      .rn_cp_iu6_i0_t1_v(rn_cp_iu6_t1_i0_t1_v),
      .rn_cp_iu6_i0_t1_t(rn_cp_iu6_t1_i0_t1_t),
      .rn_cp_iu6_i0_t1_p(rn_cp_iu6_t1_i0_t1_p),
      .rn_cp_iu6_i0_t1_a(rn_cp_iu6_t1_i0_t1_a),
      .rn_cp_iu6_i0_t2_v(rn_cp_iu6_t1_i0_t2_v),
      .rn_cp_iu6_i0_t2_t(rn_cp_iu6_t1_i0_t2_t),
      .rn_cp_iu6_i0_t2_p(rn_cp_iu6_t1_i0_t2_p),
      .rn_cp_iu6_i0_t2_a(rn_cp_iu6_t1_i0_t2_a),
      .rn_cp_iu6_i0_t3_v(rn_cp_iu6_t1_i0_t3_v),
      .rn_cp_iu6_i0_t3_t(rn_cp_iu6_t1_i0_t3_t),
      .rn_cp_iu6_i0_t3_p(rn_cp_iu6_t1_i0_t3_p),
      .rn_cp_iu6_i0_t3_a(rn_cp_iu6_t1_i0_t3_a),
      .rn_cp_iu6_i0_btb_entry(rn_cp_iu6_t1_i0_btb_entry),
      .rn_cp_iu6_i0_btb_hist(rn_cp_iu6_t1_i0_btb_hist),
      .rn_cp_iu6_i0_bta_val(rn_cp_iu6_t1_i0_bta_val),
      .rn_cp_iu6_i1_vld(rn_cp_iu6_t1_i1_vld),
      .rn_cp_iu6_i1_itag(rn_cp_iu6_t1_i1_itag),
      .rn_cp_iu6_i1_ucode(rn_cp_iu6_t1_i1_ucode),
      .rn_cp_iu6_i1_fuse_nop(rn_cp_iu6_t1_i1_fuse_nop),
      .rn_cp_iu6_i1_rte_lq(rn_cp_iu6_t1_i1_rte_lq),
      .rn_cp_iu6_i1_rte_sq(rn_cp_iu6_t1_i1_rte_sq),
      .rn_cp_iu6_i1_rte_fx0(rn_cp_iu6_t1_i1_rte_fx0),
      .rn_cp_iu6_i1_rte_fx1(rn_cp_iu6_t1_i1_rte_fx1),
      .rn_cp_iu6_i1_rte_axu0(rn_cp_iu6_t1_i1_rte_axu0),
      .rn_cp_iu6_i1_rte_axu1(rn_cp_iu6_t1_i1_rte_axu1),
      .rn_cp_iu6_i1_ifar(rn_cp_iu6_t1_i1_ifar),
      .rn_cp_iu6_i1_bta(rn_cp_iu6_t1_i1_bta),
      .rn_cp_iu6_i1_isram(rn_cp_iu6_t1_i1_isram),
      .rn_cp_iu6_i1_instr(rn_cp_iu6_t1_i1_instr),
      .rn_cp_iu6_i1_valop(rn_cp_iu6_t1_i1_valop),
      .rn_cp_iu6_i1_error(rn_cp_iu6_t1_i1_error),
      .rn_cp_iu6_i1_br_pred(rn_cp_iu6_t1_i1_br_pred),
      .rn_cp_iu6_i1_bh_update(rn_cp_iu6_t1_i1_bh_update),
      .rn_cp_iu6_i1_bh0_hist(rn_cp_iu6_t1_i1_bh0_hist),
      .rn_cp_iu6_i1_bh1_hist(rn_cp_iu6_t1_i1_bh1_hist),
      .rn_cp_iu6_i1_bh2_hist(rn_cp_iu6_t1_i1_bh2_hist),
      .rn_cp_iu6_i1_gshare(rn_cp_iu6_t1_i1_gshare),
      .rn_cp_iu6_i1_ls_ptr(rn_cp_iu6_t1_i1_ls_ptr),
      .rn_cp_iu6_i1_match(rn_cp_iu6_t1_i1_match),
      .rn_cp_iu6_i1_type_fp(rn_cp_iu6_t1_i1_type_fp),
      .rn_cp_iu6_i1_type_ap(rn_cp_iu6_t1_i1_type_ap),
      .rn_cp_iu6_i1_type_spv(rn_cp_iu6_t1_i1_type_spv),
      .rn_cp_iu6_i1_type_st(rn_cp_iu6_t1_i1_type_st),
      .rn_cp_iu6_i1_async_block(rn_cp_iu6_t1_i1_async_block),
      .rn_cp_iu6_i1_np1_flush(rn_cp_iu6_t1_i1_np1_flush),
      .rn_cp_iu6_i1_t1_v(rn_cp_iu6_t1_i1_t1_v),
      .rn_cp_iu6_i1_t1_t(rn_cp_iu6_t1_i1_t1_t),
      .rn_cp_iu6_i1_t1_p(rn_cp_iu6_t1_i1_t1_p),
      .rn_cp_iu6_i1_t1_a(rn_cp_iu6_t1_i1_t1_a),
      .rn_cp_iu6_i1_t2_v(rn_cp_iu6_t1_i1_t2_v),
      .rn_cp_iu6_i1_t2_t(rn_cp_iu6_t1_i1_t2_t),
      .rn_cp_iu6_i1_t2_p(rn_cp_iu6_t1_i1_t2_p),
      .rn_cp_iu6_i1_t2_a(rn_cp_iu6_t1_i1_t2_a),
      .rn_cp_iu6_i1_t3_v(rn_cp_iu6_t1_i1_t3_v),
      .rn_cp_iu6_i1_t3_t(rn_cp_iu6_t1_i1_t3_t),
      .rn_cp_iu6_i1_t3_p(rn_cp_iu6_t1_i1_t3_p),
      .rn_cp_iu6_i1_t3_a(rn_cp_iu6_t1_i1_t3_a),
      .rn_cp_iu6_i1_btb_entry(rn_cp_iu6_t1_i1_btb_entry),
      .rn_cp_iu6_i1_btb_hist(rn_cp_iu6_t1_i1_btb_hist),
      .rn_cp_iu6_i1_bta_val(rn_cp_iu6_t1_i1_bta_val),
      .cp_rn_empty(cp_rn_empty[1]),
      .cp_async_block(cp_async_block[1]),
      .cp_rn_i0_v(cp_rn_t1_i0_v),
      .cp_rn_i0_axu_exception_val(cp_rn_t1_i0_axu_exception_val),
      .cp_rn_i0_axu_exception(cp_rn_t1_i0_axu_exception),
      .cp_rn_i0_t1_v(cp_rn_t1_i0_t1_v),
      .cp_rn_i0_t1_t(cp_rn_t1_i0_t1_t),
      .cp_rn_i0_t1_p(cp_rn_t1_i0_t1_p),
      .cp_rn_i0_t1_a(cp_rn_t1_i0_t1_a),
      .cp_rn_i0_t2_v(cp_rn_t1_i0_t2_v),
      .cp_rn_i0_t2_t(cp_rn_t1_i0_t2_t),
      .cp_rn_i0_t2_p(cp_rn_t1_i0_t2_p),
      .cp_rn_i0_t2_a(cp_rn_t1_i0_t2_a),
      .cp_rn_i0_t3_v(cp_rn_t1_i0_t3_v),
      .cp_rn_i0_t3_t(cp_rn_t1_i0_t3_t),
      .cp_rn_i0_t3_p(cp_rn_t1_i0_t3_p),
      .cp_rn_i0_t3_a(cp_rn_t1_i0_t3_a),
      .cp_rn_i1_v(cp_rn_t1_i1_v),
      .cp_rn_i1_axu_exception_val(cp_rn_t1_i1_axu_exception_val),
      .cp_rn_i1_axu_exception(cp_rn_t1_i1_axu_exception),
      .cp_rn_i1_t1_v(cp_rn_t1_i1_t1_v),
      .cp_rn_i1_t1_t(cp_rn_t1_i1_t1_t),
      .cp_rn_i1_t1_p(cp_rn_t1_i1_t1_p),
      .cp_rn_i1_t1_a(cp_rn_t1_i1_t1_a),
      .cp_rn_i1_t2_v(cp_rn_t1_i1_t2_v),
      .cp_rn_i1_t2_t(cp_rn_t1_i1_t2_t),
      .cp_rn_i1_t2_p(cp_rn_t1_i1_t2_p),
      .cp_rn_i1_t2_a(cp_rn_t1_i1_t2_a),
      .cp_rn_i1_t3_v(cp_rn_t1_i1_t3_v),
      .cp_rn_i1_t3_t(cp_rn_t1_i1_t3_t),
      .cp_rn_i1_t3_p(cp_rn_t1_i1_t3_p),
      .cp_rn_i1_t3_a(cp_rn_t1_i1_t3_a),
      .cp_bp_val(cp_bp_t1_val),
      .cp_bp_ifar(cp_bp_t1_ifar),
      .cp_bp_bh0_hist(cp_bp_t1_bh0_hist),
      .cp_bp_bh1_hist(cp_bp_t1_bh1_hist),
      .cp_bp_bh2_hist(cp_bp_t1_bh2_hist),
      .cp_bp_br_pred(cp_bp_t1_br_pred),
      .cp_bp_br_taken(cp_bp_t1_br_taken),
      .cp_bp_bh_update(cp_bp_t1_bh_update),
      .cp_bp_bcctr(cp_bp_t1_bcctr),
      .cp_bp_bclr(cp_bp_t1_bclr),
      .cp_bp_getnia(cp_bp_t1_getnia),
      .cp_bp_group(cp_bp_t1_group),
      .cp_dis_ivax(cp_dis_ivax[1]),
      .cp_bp_lk(cp_bp_t1_lk),
      .cp_bp_bh(cp_bp_t1_bh),
      .cp_bp_gshare(cp_bp_t1_gshare),
      .cp_bp_ls_ptr(cp_bp_t1_ls_ptr),
      .cp_bp_ctr(cp_bp_t1_ctr),
      .cp_bp_btb_entry(cp_bp_t1_btb_entry),
      .cp_bp_btb_hist(cp_bp_t1_btb_hist),
      .lq0_iu_execute_vld(lq0_iu_execute_vld[1]),
      .lq0_iu_itag(lq0_iu_itag),
      .lq0_iu_n_flush(lq0_iu_n_flush),
      .lq0_iu_np1_flush(lq0_iu_np1_flush),
      .lq0_iu_dacr_type(lq0_iu_dacr_type),
      .lq0_iu_dacrw(lq0_iu_dacrw),
      .lq0_iu_instr(lq0_iu_instr),
      .lq0_iu_eff_addr(lq0_iu_eff_addr),
      .lq0_iu_exception_val(lq0_iu_exception_val),
      .lq0_iu_exception(lq0_iu_exception),
      .lq0_iu_flush2ucode(lq0_iu_flush2ucode),
      .lq0_iu_flush2ucode_type(lq0_iu_flush2ucode_type),
      .lq0_iu_recirc_val(lq0_iu_recirc_val[1]),
      .lq0_iu_dear_val(lq0_iu_dear_val[1]),
      .lq1_iu_execute_vld(lq1_iu_execute_vld[1]),
      .lq1_iu_itag(lq1_iu_itag),
      .lq1_iu_n_flush(lq1_iu_n_flush),
      .lq1_iu_np1_flush(lq1_iu_np1_flush),
      .lq1_iu_exception_val(lq1_iu_exception_val),
      .lq1_iu_exception(lq1_iu_exception),
      .lq1_iu_dacr_type(lq1_iu_dacr_type),
      .lq1_iu_dacrw(lq1_iu_dacrw),
      .lq1_iu_perf_events(lq1_iu_perf_events),
      .iu_lq_i0_completed(iu_lq_i0_completed[1]),
      .iu_lq_i1_completed(iu_lq_i1_completed[1]),
      .iu_lq_i0_completed_itag(iu_lq_t1_i0_completed_itag),
      .iu_lq_i1_completed_itag(iu_lq_t1_i1_completed_itag),
      .iu_lq_recirc_val(iu_lq_recirc_val[1]),
      .br_iu_execute_vld(br_iu_execute_vld[1]),
      .br_iu_itag(br_iu_itag),
      .br_iu_bta(br_iu_bta),
      .br_iu_redirect(br_iu_redirect[1]),
      .br_iu_taken(br_iu_taken),
      .xu_iu_execute_vld(xu_iu_execute_vld[1]),
      .xu_iu_itag(xu_iu_itag),
      .xu_iu_exception_val(xu_iu_exception_val),
      .xu_iu_exception(xu_iu_exception),
      .xu_iu_mtiar(xu_iu_mtiar[1]),
      .xu_iu_bta(xu_iu_bta),
      .xu_iu_perf_events(xu_iu_perf_events),
      .xu_iu_n_flush(xu_iu_n_flush),
      .xu_iu_np1_flush(xu_iu_np1_flush),
      .xu_iu_flush2ucode(xu_iu_flush2ucode),
      .xu1_iu_execute_vld(xu1_iu_execute_vld[1]),
      .xu1_iu_itag(xu1_iu_itag),
      .axu0_iu_execute_vld(axu0_iu_execute_vld[1]),
      .axu0_iu_itag(axu0_iu_itag),
      .axu0_iu_n_flush(axu0_iu_n_flush),
      .axu0_iu_np1_flush(axu0_iu_np1_flush),
      .axu0_iu_n_np1_flush(axu0_iu_n_np1_flush),
      .axu0_iu_exception(axu0_iu_exception),
      .axu0_iu_exception_val(axu0_iu_exception_val),
      .axu0_iu_flush2ucode(axu0_iu_flush2ucode),
      .axu0_iu_flush2ucode_type(axu0_iu_flush2ucode_type),
      .axu0_iu_async_fex(axu0_iu_async_fex[1]),
      .axu1_iu_execute_vld(axu1_iu_execute_vld[1]),
      .axu1_iu_itag(axu1_iu_itag),
      .axu1_iu_n_flush(axu1_iu_n_flush),
      .axu1_iu_np1_flush(axu1_iu_np1_flush),
      .axu1_iu_exception(axu1_iu_exception),
      .axu1_iu_exception_val(axu1_iu_exception_val),
      .axu1_iu_flush2ucode(axu1_iu_flush2ucode),
      .axu1_iu_flush2ucode_type(axu1_iu_flush2ucode_type),
      .an_ac_uncond_dbg_event(an_ac_uncond_dbg_event[1]),
      .xu_iu_external_mchk(xu_iu_external_mchk[1]),
      .xu_iu_ext_interrupt(xu_iu_ext_interrupt[1]),
      .xu_iu_dec_interrupt(xu_iu_dec_interrupt[1]),
      .xu_iu_udec_interrupt(xu_iu_udec_interrupt[1]),
      .xu_iu_perf_interrupt(xu_iu_perf_interrupt[1]),
      .xu_iu_fit_interrupt(xu_iu_fit_interrupt[1]),
      .xu_iu_crit_interrupt(xu_iu_crit_interrupt[1]),
      .xu_iu_wdog_interrupt(xu_iu_wdog_interrupt[1]),
      .xu_iu_gwdog_interrupt(xu_iu_gwdog_interrupt[1]),
      .xu_iu_gfit_interrupt(xu_iu_gfit_interrupt[1]),
      .xu_iu_gdec_interrupt(xu_iu_gdec_interrupt[1]),
      .xu_iu_dbell_interrupt(xu_iu_dbell_interrupt[1]),
      .xu_iu_cdbell_interrupt(xu_iu_cdbell_interrupt[1]),
      .xu_iu_gdbell_interrupt(xu_iu_gdbell_interrupt[1]),
      .xu_iu_gcdbell_interrupt(xu_iu_gcdbell_interrupt[1]),
      .xu_iu_gmcdbell_interrupt(xu_iu_gmcdbell_interrupt[1]),
      .xu_iu_dbsr_ide(xu_iu_dbsr_ide[1]),
      .xu_iu_rest_ifar(xu_iu_t1_rest_ifar),
      .cp_is_isync(cp_is_isync_int[1]),
      .cp_is_csync(cp_is_csync_int[1]),
      .iu_flush(iu_flush[1]),
      .cp_flush_into_uc(cp_flush_into_uc[1]),
      .cp_uc_flush_ifar(cp_uc_t1_flush_ifar),
      .cp_uc_np1_flush(cp_uc_np1_flush[1]),
      .cp_flush(cp_flush[1]),
      .cp_next_itag(cp_t1_next_itag),
      .cp_flush_itag(cp_t1_flush_itag),
      .cp_flush_ifar(cp_t1_flush_ifar),
      .cp_iu0_flush_2ucode(cp_iu0_flush_2ucode[1]),
      .cp_iu0_flush_2ucode_type(cp_iu0_flush_2ucode_type[1]),
      .cp_iu0_flush_nonspec(cp_iu0_flush_nonspec[1]),
      .pc_iu_init_reset(pc_iu_init_reset),
      .cp_rn_uc_credit_free(cp_rn_uc_credit_free[1]),
      .iu_xu_rfi(iu_xu_rfi[1]),
      .iu_xu_rfgi(iu_xu_rfgi[1]),
      .iu_xu_rfci(iu_xu_rfci[1]),
      .iu_xu_rfmci(iu_xu_rfmci[1]),
      .iu_xu_int(iu_xu_int[1]),
      .iu_xu_gint(iu_xu_gint[1]),
      .iu_xu_cint(iu_xu_cint[1]),
      .iu_xu_mcint(iu_xu_mcint[1]),
      .iu_xu_nia(iu_xu_t1_nia),
      .iu_xu_esr(iu_xu_t1_esr),
      .iu_xu_mcsr(iu_xu_t1_mcsr),
      .iu_xu_dbsr(iu_xu_t1_dbsr),
      .iu_xu_dear_update(iu_xu_dear_update[1]),
      .iu_xu_dear(iu_xu_t1_dear),
      .iu_xu_dbsr_update(iu_xu_dbsr_update[1]),
      .iu_xu_dbsr_ude(iu_xu_dbsr_ude[1]),
      .iu_xu_dbsr_ide(iu_xu_dbsr_ide[1]),
      .iu_xu_esr_update(iu_xu_esr_update[1]),
      .iu_xu_act(iu_xu_act[1]),
      .iu_xu_dbell_taken(iu_xu_dbell_taken[1]),
      .iu_xu_cdbell_taken(iu_xu_cdbell_taken[1]),
      .iu_xu_gdbell_taken(iu_xu_gdbell_taken[1]),
      .iu_xu_gcdbell_taken(iu_xu_gcdbell_taken[1]),
      .iu_xu_gmcdbell_taken(iu_xu_gmcdbell_taken[1]),
      .iu_xu_instr_cpl(iu_xu_instr_cpl[1]),
      .xu_iu_np1_async_flush(xu_iu_np1_async_flush[1]),
      .iu_xu_async_complete(iu_xu_async_complete[1]),
      .dp_cp_hold_req(dp_cp_hold_req[1]),
      .iu_mm_hold_ack(iu_mm_hold_ack[1]),
      .dp_cp_bus_snoop_hold_req(dp_cp_bus_snoop_hold_req[1]),
      .iu_mm_bus_snoop_hold_ack(iu_mm_bus_snoop_hold_ack[1]),
      .iu_spr_eheir_update(iu_spr_eheir_update[1]),
      .iu_spr_eheir(iu_spr_t1_eheir),
      .xu_iu_msr_de(xu_iu_msr_de[1]),
      .xu_iu_msr_pr(xu_iu_msr_pr[1]),
      .xu_iu_msr_cm(xu_iu_msr_cm[1]),
      .xu_iu_msr_gs(xu_iu_msr_gs[1]),
      .xu_iu_msr_me(xu_iu_msr_me[1]),
      .xu_iu_dbcr0_edm(xu_iu_dbcr0_edm[1]),
      .xu_iu_dbcr0_idm(xu_iu_dbcr0_idm[1]),
      .xu_iu_dbcr0_icmp(xu_iu_dbcr0_icmp[1]),
      .xu_iu_dbcr0_brt(xu_iu_dbcr0_brt[1]),
      .xu_iu_dbcr0_irpt(xu_iu_dbcr0_irpt[1]),
      .xu_iu_dbcr0_trap(xu_iu_dbcr0_trap[1]),
      .xu_iu_iac1_en(xu_iu_iac1_en[1]),
      .xu_iu_iac2_en(xu_iu_iac2_en[1]),
      .xu_iu_iac3_en(xu_iu_iac3_en[1]),
      .xu_iu_iac4_en(xu_iu_iac4_en[1]),
      .xu_iu_dbcr0_dac1(xu_iu_t1_dbcr0_dac1),
      .xu_iu_dbcr0_dac2(xu_iu_t1_dbcr0_dac2),
      .xu_iu_dbcr0_dac3(xu_iu_t1_dbcr0_dac3),
      .xu_iu_dbcr0_dac4(xu_iu_t1_dbcr0_dac4),
      .xu_iu_dbcr0_ret(xu_iu_dbcr0_ret[1]),
      .xu_iu_dbcr1_iac12m(xu_iu_dbcr1_iac12m[1]),
      .xu_iu_dbcr1_iac34m(xu_iu_dbcr1_iac34m[1]),
      .lq_iu_spr_dbcr3_ivc(lq_iu_spr_dbcr3_ivc[1]),
      .xu_iu_epcr_extgs(xu_iu_epcr_extgs[1]),
      .xu_iu_epcr_dtlbgs(xu_iu_epcr_dtlbgs[1]),
      .xu_iu_epcr_itlbgs(xu_iu_epcr_itlbgs[1]),
      .xu_iu_epcr_dsigs(xu_iu_epcr_dsigs[1]),
      .xu_iu_epcr_isigs(xu_iu_epcr_isigs[1]),
      .xu_iu_epcr_duvd(xu_iu_epcr_duvd[1]),
      .xu_iu_epcr_icm(xu_iu_epcr_icm[1]),
      .xu_iu_epcr_gicm(xu_iu_epcr_gicm[1]),
      .xu_iu_ccr2_en_dcr(xu_iu_spr_ccr2_en_dcr),
      .xu_iu_ccr2_ucode_dis(xu_iu_spr_ccr2_ucode_dis),
      .xu_iu_hid_mmu_mode(xu_iu_hid_mmu_mode),
      .xu_iu_xucr4_mmu_mchk(xu_iu_xucr4_mmu_mchk),
      .iu_xu_quiesce(iu_xu_quiesce[1]),
      .iu_pc_quiesce(iu_pc_quiesce[1]),
      .mm_iu_ierat_rel_val(mm_iu_ierat_rel_val[1]),
      .mm_iu_ierat_pt_fault(mm_iu_ierat_pt_fault[1]),
      .mm_iu_ierat_lrat_miss(mm_iu_ierat_lrat_miss[1]),
      .mm_iu_ierat_tlb_inelig(mm_iu_ierat_tlb_inelig[1]),
      .mm_iu_tlb_multihit_err(mm_iu_tlb_multihit_err[1]),
      .mm_iu_tlb_par_err(mm_iu_tlb_par_err[1]),
      .mm_iu_lru_par_err(mm_iu_lru_par_err[1]),
      .mm_iu_tlb_miss(mm_iu_tlb_miss[1]),
      .mm_iu_reload_hit(mm_iu_reload_hit[1]),
      .mm_iu_ierat_mmucr1(mm_iu_ierat_mmucr1[3:4]),
      .ic_cp_nonspec_hit(ic_cp_nonspec_hit[1]),
      .cp_mm_except_taken(cp_mm_except_taken_t1),
      .xu_iu_single_instr_mode(xu_iu_single_instr_mode[1]),
      .spr_single_issue(spr_single_issue[1]),
      .spr_ivpr(spr_ivpr),
      .spr_givpr(spr_givpr),
      .spr_iac1(spr_iac1),
      .spr_iac2(spr_iac2),
      .spr_iac3(spr_iac3),
      .spr_iac4(spr_iac4),
      .iu_rf_xer_p(iu_rf_t1_xer_p),
      .pc_iu_ram_active(pc_iu_ram_active[1]),
      .pc_iu_ram_flush_thread(pc_iu_ram_flush_thread[1]),
      .xu_iu_msrovride_enab(xu_iu_msrovride_enab[1]),
      .iu_pc_ram_done(iu_pc_ram_done_int[1]),
      .iu_pc_ram_interrupt(iu_pc_ram_interrupt_int[1]),
      .iu_pc_ram_unsupported(iu_pc_ram_unsupported_int[1]),
      .pc_iu_stop(pc_iu_stop[1]),
      .pc_iu_step(pc_iu_step[1]),
      .pc_iu_dbg_action(pc_iu_t1_dbg_action),
      .iu_pc_step_done(iu_pc_step_done[1]),
      .iu_pc_stop_dbg_event(iu_pc_stop_dbg_event_int[1]),
      .iu_pc_err_debug_event(iu_pc_err_debug_event[1]),
      .iu_pc_attention_instr(iu_pc_attention_instr[1]),
      .iu_pc_err_mchk_disabled(iu_pc_err_mchk_disabled[1]),
      .ac_an_debug_trigger(ac_an_debug_trigger[1]),
      .iu_xu_stop(iu_xu_stop[1])
   );
`endif


iuq_dbg iuq_cpl_dbg(
      .vdd(vdd),
      .gnd(gnd),
      .nclk(nclk),
      .thold_2(pc_iu_func_sl_thold_2),
      .pc_iu_sg_2(pc_iu_sg_2),
      .clkoff_b(clkoff_b),
      .act_dis(act_dis),
      .tc_ac_ccflush_dc(tc_ac_ccflush_dc),
      .d_mode(d_mode),
      .delay_lclkr(delay_lclkr),
      .mpw1_b(mpw1_b),
      .mpw2_b(mpw2_b),
      .func_scan_in(cp_scan_in[`THREADS]),
      .func_scan_out(cp_scan_out[`THREADS]),
      .unit_dbg_data0(unit_dbg_data0),
      .unit_dbg_data1(unit_dbg_data1),
      .unit_dbg_data2(unit_dbg_data2),
      .unit_dbg_data3(unit_dbg_data3),
      .unit_dbg_data4(unit_dbg_data4),
      .unit_dbg_data5(unit_dbg_data5),
      .unit_dbg_data6(unit_dbg_data6),
      .unit_dbg_data7(unit_dbg_data7),
      .unit_dbg_data8(unit_dbg_data8),
      .unit_dbg_data9(unit_dbg_data9),
      .unit_dbg_data10(unit_dbg_data10),
      .unit_dbg_data11(unit_dbg_data11),
      .unit_dbg_data12(unit_dbg_data12),
      .unit_dbg_data13(unit_dbg_data13),
      .unit_dbg_data14(unit_dbg_data14),
      .unit_dbg_data15(unit_dbg_data15),
      .pc_iu_trace_bus_enable(pc_iu_trace_bus_enable),
      .pc_iu_debug_mux_ctrls(pc_iu_debug_mux_ctrls),
      .debug_bus_in(debug_bus_in),
      .debug_bus_out(debug_bus_out),
      .coretrace_ctrls_in(coretrace_ctrls_in),
      .coretrace_ctrls_out(coretrace_ctrls_out)
);


endmodule
