// © IBM Corp. 2020
// This softcore is licensed under and subject to the terms of the CC-BY 4.0
// license (https://creativecommons.org/licenses/by/4.0/legalcode). 
// Additional rights, including the right to physically implement a softcore 
// that is compliant with the required sections of the Power ISA 
// Specification, will be available at no cost via the OpenPOWER Foundation. 
// This README will be updated with additional information when OpenPOWER's 
// license is available.




`include "tri_a2o.vh"




module iuq_uc_rom_even(
   vdd,
   gnd,
   nclk,
   pc_iu_func_sl_thold_0_b,
   pc_iu_sg_0,
   force_t,
   d_mode,
   delay_lclkr,
   mpw1_b,
   mpw2_b,
   scan_in,
   scan_out,
   rom_act,
   rom_addr,
   rom_data
);

    
   inout                    vdd;
    
   inout                    gnd;
    
    (* pin_data ="PIN_FUNCTION=/G_CLK/" *)
   input [0:`NCLK_WIDTH-1]  nclk;
   input                    pc_iu_func_sl_thold_0_b;
   input                    pc_iu_sg_0;
   input                    force_t;
   input                    d_mode;
   input                    delay_lclkr;
   input                    mpw1_b;
   input                    mpw2_b;
   input                    scan_in;
   output                   scan_out;

   input                    rom_act;
   input [0:9]              rom_addr;
   output [0:71]            rom_data;

   wire [1:225]             rom_instr_pt;
   wire [0:2]               count_src;
   wire                     cr_bf2fxm;
   wire                     ep;
   wire                     ext_rt;
   wire                     ext_s1;
   wire                     ext_s2;
   wire                     ext_s3;
   wire [0:9]               loop_addr;
   wire                     loop_begin;
   wire                     loop_end;
   wire [0:2]               loop_init;
   wire                     sel0_5;
   wire [0:1]               sel11_15;
   wire [0:1]               sel16_20;
   wire [0:1]               sel21_25;
   wire                     sel26_30;
   wire                     sel31;
   wire [0:1]               sel6_10;
   wire                     skip_cond;
   wire                     skip_nop;
   wire                     skip_zero;
   wire [0:31]              template;
   wire                     ucode_end;
   wire                     ucode_end_early;

   parameter                rom_addr_offset = 0;
   parameter                scan_right = rom_addr_offset + 10 - 1;

   wire [0:9]               rom_addr_d;
   wire [0:9]               rom_addr_l2;
   wire [0:scan_right]      siv;
   wire [0:scan_right]      sov;


/*
?TABLE rom_instr LISTING(final) OPTIMIZE PARMS(ON-SET, OFF-SET);
*INPUTS*========*OUTPUTS*===============================================================================================*
|               |                                                                                                       |
| rom_addr_l2   | template                         ucode_end                                                            |
| |             | |                                | ucode_end_early                                                    |
| |             | |                                | | loop_begin                                                       |
| |             | |                                | | | loop_end                                                       |
| |             | |                                | | | | count_src                                                    | -- Can DC if not (loop_begin or loop_end)
| |             | |                                | | | | |                                                            |
| |             | |                                | | | | |    ext_rt                                                  |
| |             | |                                | | | | |    | ext_s1                                                |
| |             | |                                | | | | |    | | ext_s2                                              |
| |             | |                                | | | | |    | | | ext_s3                                            |
| |             | |                                | | | | |    | | | |                                                 |
| |             | |                                | | | | |    | | | |  sel0_5                                         |
| |             | |                                | | | | |    | | | |  | sel6_10                                      |
| |             | |                                | | | | |    | | | |  | |  sel11_15                                  |
| |             | |                                | | | | |    | | | |  | |  |  sel16_20                               |
| |             | |                                | | | | |    | | | |  | |  |  |  sel21_25                            |
| |             | |                                | | | | |    | | | |  | |  |  |  |  sel26_30                         |
| |             | |                                | | | | |    | | | |  | |  |  |  |  | sel31                          |
| |             | |                                | | | | |    | | | |  | |  |  |  |  | |                              |
| |             | |                                | | | | |    | | | |  | |  |  |  |  | |  cr_bf2fxm                   |
| |             | |                                | | | | |    | | | |  | |  |  |  |  | |  | skip_cond                 |
| |             | |                                | | | | |    | | | |  | |  |  |  |  | |  | | skip_zero               | -- Can DC if loop_begin not set
| |             | |                                | | | | |    | | | |  | |  |  |  |  | |  | | | skip_nop              | -- Optimize to only be in odd side
| |             | |                                | | | | |    | | | |  | |  |  |  |  | |  | | | | loop_addr           | -- Can DC if loop_end not set; always odd side
| |             | |                                | | | | |    | | | |  | |  |  |  |  | |  | | | | |          loop_init| -- 1 less than # of times to loop; Can DC if not loop_begin or not count_src=111
| |             | |                                | | | | |    | | | |  | |  |  |  |  | |  | | | | |          |   ep   |
| |             | |         1111111111222222222233 | | | | |    | | | |  | |  |  |  |  | |  | | | | |          |   |    |
| 0123456789    | 01234567890123456789012345678901 | | | | 012  | | | |  | 01 01 01 01 | |  | | | | 0123456789 012 |    |
*TYPE*==========+=======================================================================================================+
| PPPPPPPPPP    | SSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSS S S S S SSS  S S S S  S SS SS SS SS S S  S S S S SSSSSSSSSS SSS S    |
*OPTIMIZE*----->| AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA B B B B CCC  X X X X  X XX XX XX XX X X  X X X X XXXXXXXXXX XYX X    |
*TERMS*=========+=======================================================================================================+
| 0000000000    | 00111000000--------------------- 0 0 0 - ---  1 0 - -  0 00 01 01 01 1 1  0 0 - 0 ---------- --- -    | # addi s0,RA,D 	-lhz,lhzu
| 0000000010    | 10001000010000000000000000000001 0 0 0 - ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # lbz s2,1(s0)
| 0000000100    | 01010100010000100100010000101110 0 0 0 - ---  1 1 - -  0 00 00 00 00 0 0  0 1 - 0 ---------- --- -    | # rlwinm s2,s2,8,16,23 	-skip_c
| 0000000110    | 01101000010-----0000000000000000 0 1 0 - ---  0 1 - -  0 00 11 00 00 0 0  0 0 - 0 ---------- --- -    | # xori RT,s2,0 	-end for non-update

| 0000010000    | 011111-----00000-----00000111000 0 0 0 - ---  1 0 0 -  0 11 00 01 00 0 0  0 0 - 0 ---------- --- 0    | # and s0,RB,RB 	-lhzx,lhzux,lhbrx
| 0000010010    | 00111000011000000000000000000001 0 0 0 - ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- 0    | # addi s3,s0,1
| 0000010100    | 01010000001000100100010000101110 0 0 0 - ---  1 1 1 -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- 0    | # rlwimi s2,s1,8,16,23
| 0000010110    | 01111100010000100000101101111000 0 0 0 - ---  1 1 1 -  0 00 00 00 00 0 0  0 1 - 0 ---------- --- 0    | # or s2,s2,s1 	-skip_c
| 0000011000    | 011111----------0000001000010100 1 - 0 - ---  0 0 1 -  0 10 01 00 00 0 0  0 0 - 0 ---------- --- 0    | # add RA,RA,s0

| 0000100000    | 00111000000--------------------- 0 0 0 - ---  1 0 - -  0 00 01 01 01 1 1  0 0 - 0 ---------- --- -    | # addi s0,RA,D 	-lha,lhau
| 0000100010    | 10001000010000000000000000000001 0 0 0 - ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # lbz s2,1(s0)
| 0000100100    | 01010100010000100100010000101110 0 0 0 - ---  1 1 - -  0 00 00 00 00 0 0  0 1 - 0 ---------- --- -    | # rlwinm s2,s2,8,16,23 	-skip_c
| 0000100110    | 01111100010----------11100110100 0 1 0 - ---  0 1 - -  0 00 11 -- 00 0 0  0 0 - 0 ---------- --- -    | # extsh RT,s2 	-end for non-update

| 0000110000    | 00111000000-----0000000000000000 0 0 0 - ---  1 0 - -  0 00 01 00 00 0 0  0 0 - 0 ---------- --- -    | # addi s0,RA,0 	-lhax,lhaux
| 0000110010    | 10001000001000000000000000000000 0 0 0 - ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # lbz s1,0(s0)
| 0000110100    | 01010000001000100100010000101110 0 0 0 - ---  1 1 1 -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # rlwimi s2,s1,8,16,23
| 0000110110    | 01111100010000100000101101111000 0 0 0 - ---  1 1 1 -  0 00 00 00 00 0 0  0 1 - 0 ---------- --- -    | # or s2,s2,s1 	-skip_c
| 0000111000    | 01101000000-----0000000000000000 1 - 0 - ---  0 1 - -  0 00 01 00 00 0 0  0 0 - 0 ---------- --- -    | # xori RA,s0,0

| 0001000000    | 00111000000--------------------- 0 0 0 - ---  1 0 - -  0 00 01 01 01 1 1  0 0 - 0 ---------- --- -    | # addi s0,RA,D 	-lwz,lwzu
| 0001000010    | 00111000000000000000000000000001 0 0 1 0 111  1 1 - -  0 00 00 00 00 0 0  0 0 0 0 ---------- 010 -    | # addi s0,s0,1 	-loop_begin,cnt=3
| 0001000100    | 10001000001000000000000000000000 0 0 0 0 ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # lbz s1,0(s0)
| 0001000110    | 01010100010000100100000000111110 0 0 0 - ---  1 1 - -  0 00 00 00 00 0 0  0 1 - 0 ---------- --- -    | # rlwinm s2,s2,8,0,31 	-skip_c
| 0001001000    | 01010000001000101100000000001110 0 0 0 - ---  1 1 1 -  0 00 00 00 00 0 0  0 1 - 0 ---------- --- -    | # rlwimi s2,s1,24,0,7 	-skip_c
| 0001001010    | 001110-------------------------- 1 - 0 - ---  0 0 - -  0 10 01 01 01 1 1  0 0 - 0 ---------- --- -    | # addi RA,RA,D

| 0001010000    | 011111-----00000-----00000111000 0 0 0 - ---  1 0 0 -  0 11 00 01 00 0 0  0 0 - 0 ---------- --- 0    | # and s0,RB,RB 	-lwzx,lwzux,lwbrx
| 0001010010    | 00111000000000000000000000000001 0 0 1 0 111  1 1 - -  0 00 00 00 00 0 0  0 0 0 0 ---------- 010 0    | # addi s0,s0,1 	-loop_begin,cnt=3
| 0001010100    | 01111100001-----000000001010111- 0 0 0 0 ---  1 0 1 -  0 00 01 00 00 0 -  0 0 - 0 ---------- --- 1    | # lbzx s1,RA,s0
| 0001010110    | 01010100010000100100000000111110 0 0 0 - ---  1 1 - -  0 00 00 00 00 0 0  0 1 - 0 ---------- --- 0    | # rlwinm s2,s2,8,0,31 	-skip_c
| 0001011000    | 01010000001000101100000000001110 0 0 0 - ---  1 1 1 -  0 00 00 00 00 0 0  0 1 - 0 ---------- --- 0    | # rlwimi s2,s1,24,0,7 	-skip_c
| 0001011010    | 00111000001-----1111111111111101 0 - 0 - ---  1 0 - -  0 00 01 00 00 0 0  0 0 - 0 ---------- --- 0    | # addi s1,RA,-3

| 0001100000    | 00111000000-----1111111111111110 0 - 0 - ---  1 0 - -  0 00 01 00 00 0 0  0 0 - 0 ---------- --- -    | # addi s0,RA,-2 	-lwa
| 0001100010    | 00111000000000000000000000000001 0 - 1 0 111  1 1 - -  0 00 00 00 00 0 0  0 0 0 0 ---------- 010 -    | # addi s0,s0,1 	-loop_begin,cnt=3
| 0001100100    | 1000100000100000---------------- 0 - 0 0 ---  1 1 - -  0 00 00 01 01 1 1  0 0 - 0 ---------- --- -    | # lbz s1,D(s0)
| 0001100110    | 01010100010000100100000000111110 0 - 0 - ---  1 1 - -  0 00 00 00 00 0 0  0 1 - 0 ---------- --- -    | # rlwinm s2,s2,8,0,31 	-skip_c
| 0001101000    | 01010000001000101100000000001110 0 - 0 - ---  1 1 1 -  0 00 00 00 00 0 0  0 1 - 0 ---------- --- -    | # rlwimi s2,s1,24,0,7 	-skip_c

| 0001110000    | 011111-----00000-----00000111000 0 0 0 - ---  1 0 0 -  0 11 00 01 00 0 0  0 0 - 0 ---------- --- -    | # and s0,RB,RB 	-lwax,lwaux
| 0001110010    | 00111000000000000000000000000001 0 0 1 0 111  1 1 - -  0 00 00 00 00 0 0  0 0 0 0 ---------- 010 -    | # addi s0,s0,1 	-loop_begin,cnt=3
| 0001110100    | 01111100001-----000000001010111- 0 0 0 0 ---  1 0 1 -  0 00 01 00 00 0 -  0 0 - 0 ---------- --- -    | # lbzx s1,RA,s0
| 0001110110    | 01010100010000100100000000111110 0 0 0 - ---  1 1 - -  0 00 00 00 00 0 0  0 1 - 0 ---------- --- -    | # rlwinm s2,s2,8,0,31 	-skip_c
| 0001111000    | 01010000001000101100000000001110 0 0 0 - ---  1 1 1 -  0 00 00 00 00 0 0  0 1 - 0 ---------- --- -    | # rlwimi s2,s1,24,0,7 	-skip_c
| 0001111010    | 00111000001-----1111111111111101 0 - 0 - ---  1 0 - -  0 00 01 00 00 0 0  0 0 - 0 ---------- --- -    | # addi s1,RA,-3

| 0010000000    | 00111000000--------------------0 0 0 0 - ---  1 0 - -  0 00 01 01 01 1 0  0 0 - 0 ---------- --- -    | # addi s0,RA,DS 	-ld,ldu
| 0010000010    | 00111000000000000000000000000001 0 0 1 0 111  1 1 - -  0 00 00 00 00 0 0  0 0 0 0 ---------- 110 -    | # addi s0,s0,1 	-loop_begin,cnt=7
| 0010000100    | 10001000001000000000000000000000 0 0 0 0 ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # lbz s1,0(s0)
| 0010000110    | 01111000010000101100000000000010 0 0 1 0 111  1 1 - -  0 00 00 00 00 0 0  0 1 0 0 ---------- 110 -    | # rldicl s2,s2,56,0 	-skip_c,loop_begin,cnt=7
| 0010001000    | 01010000010000010000011000111110 0 0 0 1 ---  1 1 1 -  0 00 00 00 00 0 0  0 1 - 0 ---------- --- -    | # rlwimi s1,s2,0,24,31 	-skip_c,loop_end
| 0010001010    | 01101000010-----0000000000000000 0 1 0 - ---  0 1 - -  0 00 11 00 00 0 0  0 0 - 0 ---------- --- -    | # xori RT,s2,0 	-end for non-update

| 0010010000    | 011111-----00000-----00000111000 0 0 0 - ---  1 0 0 -  0 11 00 01 00 0 0  0 0 - 0 ---------- --- 0    | # and s0,RB,RB 	-ldx,ldux,ldbrx
| 0010010010    | 00111000000000000000000000000001 0 0 1 0 111  1 1 - -  0 00 00 00 00 0 0  0 0 0 0 ---------- 110 0    | # addi s0,s0,1 	-loop_begin,cnt=7
| 0010010100    | 01111100001-----000000001010111- 0 0 0 0 ---  1 0 1 -  0 00 01 00 00 0 -  0 0 - 0 ---------- --- 1    | # lbzx s1,RA,s0
| 0010010110    | 01111000010000101100000000000010 0 0 1 0 111  1 1 - -  0 00 00 00 00 0 0  0 1 0 0 ---------- 110 0    | # rldicl s2,s2,56,0 	-skip_c,loop_begin,cnt=7
| 0010011000    | 01010000010000010000011000111110 0 0 0 1 ---  1 1 1 -  0 00 00 00 00 0 0  0 1 - 0 ---------- --- 0    | # rlwimi s1,s2,0,24,31 	-skip_c,loop_end
| 0010011010    | 01101000010-----0000000000000000 0 1 0 - ---  0 1 - -  0 00 11 00 00 0 0  0 0 - 0 ---------- --- 0    | # xori RT,s2,0 	-end for non-update
| 0010011100    | 011111-----000010000001000010100 1 - 0 - ---  0 1 1 -  0 10 00 00 00 0 0  0 0 - 0 ---------- --- 0    | # add RA,s1,s0

| 0010100000    | 00111000000--------------------- 0 - 0 - ---  1 0 - -  0 00 01 01 01 1 1  0 0 - 0 ---------- --- -    | # addi s0,RA,D 	-lmw
| 0010100010    | 100000-----000000000000000000000 0 - 1 0 100  0 1 - -  0 01 00 00 00 0 0  0 0 1 0 ---------- --- -    | # lwz RT,0(s0) 	-loop_begin,skip_zero
| 0010100100    | 100000-----000000000000000000000 1 - 0 - ---  0 1 - -  0 01 00 00 00 0 0  0 0 - 0 ---------- --- -    | # lwz RT,0(s0)

| 0010110000    | 00111000000-----0000000000000000 0 - 0 - ---  1 0 - -  0 00 01 00 00 0 0  0 0 - 0 ---------- --- -    | # addi s0,RA,0 	-lswi
| 0010110010    | 10001000010000000000000000000000 0 - 1 0 101  1 1 - -  0 00 00 00 00 0 0  0 0 1 0 ---------- --- -    | # lbz s2,0(s0) 	-loop_begin,skip_zero
| 0010110100    | 10001000001000000000000000000001 0 - 0 0 ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # lbz s1,1(s0)
| 0010110110    | 10001000001000000000000000000010 0 - 0 0 ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # lbz s1,2(s0)
| 0010111000    | 10001000001000000000000000000011 0 - 0 0 ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # lbz s1,3(s0)
| 0010111010    | 01111100010-----0000101101111000 0 - 0 1 ---  0 1 1 -  0 00 11 00 00 0 0  0 0 - 0 ---------- --- -    | # or RT,s2,s1 	-loop_end
| 0010111100    | 10001000001000000000000000000000 0 - 1 0 000  1 1 - -  0 00 00 00 00 0 0  0 0 0 0 ---------- --- -    | # lbz s1,0(s0) 	-loop_begin
| 0010111110    | 00111000000000000000000000000001 0 - 0 0 ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # addi s0,s0,1
| 0011000000    | 01010100010000100100000000101110 0 - 1 0 001  1 1 - -  0 00 00 00 00 0 0  0 0 1 0 ---------- --- -    | # rlwinm s2,s2,8,0,23 	-loop_begin,skip_zero
| 0011000010    | 01101000010-----0000000000000000 1 - 0 - ---  0 1 - -  0 00 11 00 00 0 0  0 0 - 0 ---------- --- -    | # xori RT,s2,0

| 0011010000    | 00111000010000000000000000000000 0 - 0 - ---  1 0 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # addi s2,R0,0 	-lswx
| 0011010010    | 0111110001000000-----0001010111- 0 - 1 0 110  1 1 0 -  0 00 00 01 00 0 -  0 0 1 0 ---------- --- -    | # lbzx s2,s0,RB 	-loop_begin,skip_zero
| 0011010100    | 01010100010000101100000000111110 0 - 0 0 ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # rlwinm s2,s2,24,0,31
| 0011010110    | 00111000000000000000000000000001 0 - 0 0 ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # addi s0,s0,1
| 0011011000    | 0111110000100000-----0001010111- 0 - 0 0 ---  1 1 0 -  0 00 00 01 00 0 -  0 0 - 0 ---------- --- -    | # lbzx s1,s0,RB
| 0011011010    | 01010000001000100100010000101110 0 - 0 0 ---  1 1 1 -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # rlwimi s2,s1,8,16,23
| 0011011100    | 00111000000000000000000000000001 0 - 0 0 ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # addi s0,s0,1
| 0011011110    | 0111110000100000-----0001010111- 0 - 1 0 010  1 1 0 -  0 00 00 01 00 0 -  0 0 1 0 ---------- --- -    | # lbzx s1,s0,RB 	-loop_begin,skip_zero
| 0011100000    | 00111000000000000000000000000001 0 - 0 0 ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # addi s0,s0,1
| 0011100010    | 01010100010000100100000000101110 0 - 1 0 011  1 1 - -  0 00 00 00 00 0 0  0 0 1 0 ---------- --- -    | # rlwinm s2,s2,8,0,23 	-loop_begin,skip_zero
| 0011100100    | 01101000010-----0000000000000000 1 - 0 - ---  0 1 - -  0 00 11 00 00 0 0  0 0 - 0 ---------- --- -    | # xori RT,s2,0


| 0100000000    | 010101-----000101100000000111110 0 0 0 - ---  1 0 - -  0 01 00 00 00 0 0  0 0 - 0 ---------- --- -    | # rlwinm s2,RS,24,0,31 	-sth,sthu
| 0100000010    | 010101-----000101000000000001110 0 0 0 - ---  1 0 - -  0 01 00 00 00 0 0  0 1 - 0 ---------- --- -    | # rlwinm s2,RS,16,0,7 	-skip_c
| 0100000100    | 10011000010000000000000000000000 0 0 0 - ---  - 1 - 1  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # stb s2,0(s0)
| 0100000110    | 10011000010000000000000000000001 0 1 0 - ---  - 1 - 1  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # stb s2,1(s0) 	-end for non-update

| 0100010000    | 010101-----000101100000000111110 0 0 0 - ---  1 0 - -  0 01 00 00 00 0 0  0 0 - 0 ---------- --- 0    | # rlwinm s2,RS,24,0,31 	-sthx,sthux,sthbrx
| 0100010010    | 010101-----000101000000000001110 0 0 0 - ---  1 0 - -  0 01 00 00 00 0 0  0 1 - 0 ---------- --- 0    | # rlwinm s2,RS,16,0,7 	-skip_c
| 0100010100    | 01111100010----------0011010111- 0 0 0 - ---  - 0 0 1  0 00 01 01 00 0 -  0 0 - 0 ---------- --- 1    | # stbx s2,RA,RB
| 0100010110    | 0111110001000000-----0011010111- 0 1 0 - ---  - 1 0 1  0 00 00 01 00 0 -  0 0 - 0 ---------- --- 1    | # stbx s2,s0,RB 	-end for non-update
| 0100011000    | 011111-----00000-----01000010100 1 - 0 - ---  0 1 0 -  0 10 00 01 00 0 0  0 0 - 0 ---------- --- 0    | # add RA,s0,RB

| 0101000000    | 010101-----000100100000000111110 0 0 0 - ---  1 0 - -  0 01 00 00 00 0 0  0 0 - 0 ---------- --- -    | # rlwinm s2,RS,8,0,31 	-stw,stwu
| 0101000010    | 01010000010000101000010000101110 0 0 0 - ---  1 1 1 -  0 00 00 00 00 0 0  0 1 - 0 ---------- --- -    | # rlwimi s2,s2,16,16,23 	-skip_c
| 0101000100    | 00111000000--------------------- 0 0 0 - ---  1 0 - -  0 00 01 01 01 1 1  0 0 - 0 ---------- --- -    | # addi s0,RA,D
| 0101000110    | 00111000000000000000000000000001 0 0 1 0 111  1 1 - -  0 00 00 00 00 0 0  0 0 0 0 ---------- 010 -    | # addi s0,s0,1 	-loop_begin,cnt=3
| 0101001000    | 10011000010000000000000000000000 0 1 0 1 ---  - 1 - 1  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # stb s2,0(s0) 	-loop_end,end for non-update

| 0101010000    | 010101-----000100100000000111110 0 0 0 - ---  1 0 - -  0 01 00 00 00 0 0  0 0 - 0 ---------- --- 0    | # rlwinm s2,RS,8,0,31 	-stwx,stwux,stwbrx
| 0101010010    | 01010000010000101000010000101110 0 0 0 - ---  1 1 1 -  0 00 00 00 00 0 0  0 1 - 0 ---------- --- 0    | # rlwimi s2,s2,16,16,23 	-skip_c
| 0101010100    | 00111000000-----0000000000000000 0 0 0 - ---  1 0 - -  0 00 01 00 00 0 0  0 0 - 0 ---------- --- 0    | # addi s0,RA,0
| 0101010110    | 00111000000000000000000000000001 0 0 1 0 111  1 1 - -  0 00 00 00 00 0 0  0 0 0 0 ---------- 010 0    | # addi s0,s0,1 	-loop_begin,cnt=3
| 0101011000    | 0111110001000000-----0011010111- 0 1 0 1 ---  - 1 0 1  0 00 00 01 00 0 -  0 0 - 0 ---------- --- 1    | # stbx s2,s0,RB 	-loop_end,end for non-update

| 0110000000    | 011110-----000100100000000000000 0 0 0 - ---  1 0 - -  0 01 00 00 00 0 0  0 0 - 0 ---------- --- -    | # rldicl s2,RS,8,0 	-std,stdu
| 0110000010    | 01111000010000101100000000000010 0 0 1 0 111  1 1 - -  0 00 00 00 00 0 0  0 1 0 0 ---------- 111 -    | # rldicl s2,s2,56,0 	-skip_c,loop_begin,cnt=8
| 0110000100    | 01010000010000010000011000111110 0 0 0 1 ---  1 1 1 -  0 00 00 00 00 0 0  0 1 - 0 ---------- --- -    | # rlwimi s1,s2,0,24,31 	-skip_c,loop_end
| 0110000110    | 1001100001000000---------------0 0 0 1 0 111  - 1 - 1  0 00 00 01 01 1 0  0 0 0 0 ---------- 110 -    | # stb s2,DS(s0) 	-loop_begin,cnt=7
| 0110001000    | 01111000010000100100000000000000 0 0 0 1 ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # rldicl s2,s2,8,0 	-loop_end
| 0110001010    | 001110-------------------------0 1 - 0 - ---  0 0 - -  0 10 01 01 01 1 0  0 0 - 0 ---------- --- -    | # addi RA,RA,DS

| 0110010000    | 011110-----000100100000000000000 0 0 0 - ---  1 0 - -  0 01 00 00 00 0 0  0 0 - 0 ---------- --- 0    | # rldicl s2,RS,8,0 	-stdx,stdux,stdbrx
| 0110010010    | 01111000010000101100000000000010 0 0 1 0 111  1 1 - -  0 00 00 00 00 0 0  0 1 0 0 ---------- 111 0    | # rldicl s2,s2,56,0 	-skip_c,loop_begin,cnt=8
| 0110010100    | 01010000010000010000011000111110 0 0 0 1 ---  1 1 1 -  0 00 00 00 00 0 0  0 1 - 0 ---------- --- 0    | # rlwimi s1,s2,0,24,31 	-skip_c,loop_end
| 0110010110    | 0111110001000000-----0011010111- 0 0 1 0 111  - 1 0 1  0 00 00 01 00 0 -  0 0 0 0 ---------- 110 1    | # stbx s2,s0,RB 	-loop_begin,cnt=7
| 0110011000    | 01111000010000100100000000000000 0 0 0 1 ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- 0    | # rldicl s2,s2,8,0 	-loop_end
| 0110011010    | 011111---------------01000010100 1 - 0 - ---  0 0 0 -  0 10 01 01 00 0 0  0 0 - 0 ---------- --- 0    | # add RA,RA,RB


| 0110100000    | 00111000000--------------------- 0 - 0 - ---  1 0 - -  0 00 01 01 01 1 1  0 0 - 0 ---------- --- -    | # addi s0,RA,D 	-stmw
| 0110100010    | 100100-----000000000000000000000 0 - 1 0 100  - 1 - 0  0 01 00 00 00 0 0  0 0 1 0 ---------- --- -    | # stw RS,0(s0) 	-loop_begin,skip_zero
| 0110100100    | 100100-----000000000000000000000 1 - 0 - ---  - 1 - 0  0 01 00 00 00 0 0  0 0 - 0 ---------- --- -    | # stw RS,0(s0)

| 0110110000    | 00111000000-----0000000000000000 0 - 0 - ---  1 0 - -  0 00 01 00 00 0 0  0 0 - 0 ---------- --- -    | # addi s0,RA,0 	-stswi
| 0110110010    | 010101-----000100100000000111110 0 - 1 0 101  1 0 - -  0 01 00 00 00 0 0  0 0 1 0 ---------- --- -    | # rlwinm s2,RS,8,0,31 	-loop_begin,skip_zero
| 0110110100    | 01010100010000100100000000111110 0 - 0 0 ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # rlwinm s2,s2,8,0,31
| 0110110110    | 01010100010000100100000000111110 0 - 0 0 ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # rlwinm s2,s2,8,0,31
| 0110111000    | 01010100010000100100000000111110 0 - 0 0 ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # rlwinm s2,s2,8,0,31
| 0110111010    | 00111000000000000000000000000100 0 - 0 1 ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # addi s0,s0,4 	-loop_end
| 0110111100    | 010101-----000100100000000111110 0 - 0 - ---  1 0 - -  0 01 00 00 00 0 0  0 0 - 0 ---------- --- -    | # rlwinm s2,RS,8,0,31
| 0110111110    | 10011000010000000000000000000000 0 - 1 0 000  - 1 - 1  0 00 00 00 00 0 0  0 0 0 0 ---------- --- -    | # stb s2,0(s0) 	-loop_begin
| 0111000000    | 01010100010000100100000000111110 1 - 0 1 ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # rlwinm s2,s2,8,0,31 	-loop_end

| 0111010000    | 00111000000-----0000000000000000 0 - 0 - ---  1 0 - -  0 00 01 00 00 0 0  0 0 - 0 ---------- --- -    | # addi s0,RA,0 	-stswx
| 0111010010    | 010101-----000100100000000111110 0 - 1 0 110  1 0 - -  0 01 00 00 00 0 0  0 0 1 0 ---------- --- -    | # rlwinm s2,RS,8,0,31 	-loop_begin,skip_zero
| 0111010100    | 00111000000000000000000000000001 0 - 0 0 ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # addi s0,s0,1
| 0111010110    | 0111110001000000-----0011010111- 0 - 0 0 ---  - 1 0 1  0 00 00 01 00 0 -  0 0 - 0 ---------- --- -    | # stbx s2,s0,RB
| 0111011000    | 01010100010000100100000000111110 0 - 0 0 ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # rlwinm s2,s2,8,0,31
| 0111011010    | 00111000000000000000000000000001 0 - 0 0 ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # addi s0,s0,1
| 0111011100    | 0111110001000000-----0011010111- 0 - 0 0 ---  - 1 0 1  0 00 00 01 00 0 -  0 0 - 0 ---------- --- -    | # stbx s2,s0,RB
| 0111011110    | 010101-----000100100000000111110 0 - 0 - ---  1 0 - -  0 01 00 00 00 0 0  0 0 - 0 ---------- --- -    | # rlwinm s2,RS,8,0,31
| 0111100000    | 0111110001000000-----0011010111- 0 - 1 0 010  - 1 0 1  0 00 00 01 00 0 -  0 0 1 0 ---------- --- -    | # stbx s2,s0,RB 	-loop_begin,skip_zero
| 0111100010    | 01010100010000100100000000111110 0 - 0 1 ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # rlwinm s2,s2,8,0,31 	-loop_end


| 0101100000    | 0111110000000001000000101010011- 0 - 0 - ---  1 - - -  0 00 00 00 00 0 -  0 0 - 0 ---------- --- -    | # mfxer s0 	-mcrxr
| 0101100010    | 01111100000000100000101001111000 0 - 0 - ---  1 1 1 -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # xor s2,s0,s1
| 0101100100    | 01111100000000010000101101111000 0 - 0 - ---  1 1 1 -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # or s1,s0,s1
| 0101100110    | 01111100000000010000101101111000 0 - 0 - ---  1 1 1 -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # or s1,s0,s1
| 0101101000    | 01111100000000010000101101111000 0 - 0 - ---  1 1 1 -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # or s1,s0,s1
| 0101101010    | 0111110001000001000000111010011- 1 - 0 - ---  - 1 - -  0 00 00 00 00 0 -  0 0 - 0 ---------- --- -    | # mtxer s2

| 0101110000    | 011111-----110000000-0000010011- 0 - 0 - ---  0 - - -  0 01 00 00 00 0 -  0 0 - 0 ---------- --- -    | # mfocrf RT,0x80      -mfcr
| 0101110010    | 011111----------0000001101111000 0 - 0 - ---  0 0 1 -  0 01 11 00 00 0 0  0 0 - 0 ---------- --- -    | # or RT,RT,s0
| 0101110100    | 011111----------0000001101111000 0 - 0 - ---  0 0 1 -  0 01 11 00 00 0 0  0 0 - 0 ---------- --- -    | # or RT,RT,s0
| 0101110110    | 011111----------0000001101111000 0 - 0 - ---  0 0 1 -  0 01 11 00 00 0 0  0 0 - 0 ---------- --- -    | # or RT,RT,s0
| 0101111000    | 011111----------0000001101111000 0 - 0 - ---  0 0 1 -  0 01 11 00 00 0 0  0 0 - 0 ---------- --- -    | # or RT,RT,s0
| 0101111010    | 011111----------0000001101111000 0 - 0 - ---  0 0 1 -  0 01 11 00 00 0 0  0 0 - 0 ---------- --- -    | # or RT,RT,s0
| 0101111100    | 011111----------0000001101111000 0 - 0 - ---  0 0 1 -  0 01 11 00 00 0 0  0 0 - 0 ---------- --- -    | # or RT,RT,s0
| 0101111110    | 011111----------0000001101111000 1 - 0 - ---  0 0 1 -  0 01 11 00 00 0 0  0 0 - 0 ---------- --- -    | # or RT,RT,s0


| 0111110000    | 011111-----110000000-0010010000- 0 - 0 - ---  - 0 - -  0 01 00 00 00 0 -  0 0 - 0 ---------- --- -    | # mtocrf 0x80,RS      -mtcrf
| 0111110010    | 011111-----100100000-0010010000- 0 - 0 - ---  - 0 - -  0 01 00 00 00 0 -  0 0 - 0 ---------- --- -    | # mtocrf 0x20,RS
| 0111110100    | 011111-----100001000-0010010000- 0 - 0 - ---  - 0 - -  0 01 00 00 00 0 -  0 0 - 0 ---------- --- -    | # mtocrf 0x08,RS
| 0111110110    | 011111-----100000010-0010010000- 0 - 0 - ---  - 0 - -  0 01 00 00 00 0 -  0 0 - 0 ---------- --- -    | # mtocrf 0x02,RS



| 1010100000    | 100010-------------------------- 0 - 0 - ---  0 0 - -  0 01 01 01 01 1 1  0 0 - 0 ---------- --- -    | # lbz RT,D(RA) 	-lbzu

| 1010101000    | 01111100000----------01000010100 0 - 0 - ---  1 0 0 -  0 00 01 01 00 0 0  0 0 - 0 ---------- --- -    | # add s0,RA,RB 	-lbzux
| 1010101010    | 01101000000-----0000000000000000 1 - 0 - ---  0 1 - -  0 00 01 00 00 0 0  0 0 - 0 ---------- --- -    | # xori RA,s0,0

| 1010110000    | 101000-------------------------- 0 - 0 - ---  0 0 - -  0 01 01 01 01 1 1  0 0 - 0 ---------- --- -    | # lhz RT,D(RA) 	-lhzu

| 1010111000    | 01111100000----------01000010100 0 - 0 - ---  1 0 0 -  0 00 01 01 00 0 0  0 0 - 0 ---------- --- -    | # add s0,RA,RB 	-lhzux
| 1010111010    | 01101000000-----0000000000000000 1 - 0 - ---  0 1 - -  0 00 01 00 00 0 0  0 0 - 0 ---------- --- -    | # xori RA,s0,0

| 1011000000    | 100000-------------------------- 0 - 0 - ---  0 0 - -  0 01 01 01 01 1 1  0 0 - 0 ---------- --- -    | # lwz RT,D(RA) 	-lwzu

| 1011001000    | 01111100000----------01000010100 0 - 0 - ---  1 0 0 -  0 00 01 01 00 0 0  0 0 - 0 ---------- --- -    | # add s0,RA,RB 	-lwzux
| 1011001010    | 01101000000-----0000000000000000 1 - 0 - ---  0 1 - -  0 00 01 00 00 0 0  0 0 - 0 ---------- --- -    | # xori RA,s0,0

| 1011010000    | 111010-------------------------0 0 - 0 - ---  0 0 - -  0 01 01 01 01 1 0  0 0 - 0 ---------- --- -    | # ld RT,DS(RA) 	-ldu

| 1011011000    | 01111100000----------01000010100 0 - 0 - ---  1 0 0 -  0 00 01 01 00 0 0  0 0 - 0 ---------- --- -    | # add s0,RA,RB 	-ldux
| 1011011010    | 01101000000-----0000000000000000 1 - 0 - ---  0 1 - -  0 00 01 00 00 0 0  0 0 - 0 ---------- --- -    | # xori RA,s0,0

| 1011100000    | 101010-------------------------- 0 - 0 - ---  0 0 - -  0 01 01 01 01 1 1  0 0 - 0 ---------- --- -    | # lha RT,D(RA) 	-lhau

| 1011101000    | 01111100000----------01000010100 0 - 0 - ---  1 0 0 -  0 00 01 01 00 0 0  0 0 - 0 ---------- --- -    | # add s0,RA,RB 	-lhaux
| 1011101010    | 01101000000-----0000000000000000 1 - 0 - ---  0 1 - -  0 00 01 00 00 0 0  0 0 - 0 ---------- --- -    | # xori RA,s0,0

| 1011111000    | 01111100000----------01000010100 0 - 0 - ---  1 0 0 -  0 00 01 01 00 0 0  0 0 - 0 ---------- --- -    | # add s0,RA,RB 	-lwaux
| 1011111010    | 01101000000-----0000000000000000 1 - 0 - ---  0 1 - -  0 00 01 00 00 0 0  0 0 - 0 ---------- --- -    | # xori RA,s0,0



| 1000110000    | 011111-----00000-----00000111000 0 - 0 - ---  1 0 0 -  0 11 00 01 00 0 0  0 0 - 0 ---------- --- -    | # and s0,RB,RB        -lfiwax
| 1000110010    | 00111000000000000000000000000001 0 - 1 0 111  1 1 - -  0 00 00 00 00 0 0  0 0 0 0 ---------- 010 -    | # addi s0,s0,1 	-loop_begin,cnt=3
| 1000110100    | 01111100001-----000000001010111- 0 - 0 0 ---  1 0 1 -  0 00 01 00 00 0 -  0 0 - 0 ---------- --- -    | # lbzx s1,RA,s0
| 1000110110    | 01010100010000100100000000111110 0 - 0 - ---  1 1 - -  0 00 00 00 00 0 0  0 1 - 0 ---------- --- -    | # rlwinm s2,s2,8,0,31 	-skip_c
| 1000111000    | 01010000001000101100000000001110 0 - 0 - ---  1 1 1 -  0 00 00 00 00 0 0  0 1 - 0 ---------- --- -    | # rlwimi s2,s1,24,0,7 	-skip_c

| 1001110000    | 011111-----00000-----00000111000 0 - 0 - ---  1 0 0 -  0 11 00 01 00 0 0  0 0 - 0 ---------- --- -    | # and s0,RB,RB        -lfiwzx
| 1001110010    | 00111000000000000000000000000001 0 - 1 0 111  1 1 - -  0 00 00 00 00 0 0  0 0 0 0 ---------- 010 -    | # addi s0,s0,1 	-loop_begin,cnt=3
| 1001110100    | 01111100001-----000000001010111- 0 - 0 0 ---  1 0 1 -  0 00 01 00 00 0 -  0 0 - 0 ---------- --- -    | # lbzx s1,RA,s0
| 1001110110    | 01010100010000100100000000111110 0 - 0 - ---  1 1 - -  0 00 00 00 00 0 0  0 1 - 0 ---------- --- -    | # rlwinm s2,s2,8,0,31 	-skip_c
| 1001111000    | 01010000001000101100000000001110 0 - 0 - ---  1 1 1 -  0 00 00 00 00 0 0  0 1 - 0 ---------- --- -    | # rlwimi s2,s1,24,0,7 	-skip_c

| 1001000000    | 00111000000--------------------- 0 0 0 - ---  1 0 - -  0 00 01 01 01 1 1  0 0 - 0 ---------- --- -    | # addi s0,RA,D 	-lfs,lfsu
| 1001000010    | 00111000000000000000000000000001 0 0 1 0 111  1 1 - -  0 00 00 00 00 0 0  0 0 0 0 ---------- 010 -    | # addi s0,s0,1 	-loop_begin,cnt=3
| 1001000100    | 10001000001000000000000000000000 0 0 0 0 ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # lbz s1,0(s0)
| 1001000110    | 01010100010000100100000000111110 0 0 0 - ---  1 1 - -  0 00 00 00 00 0 0  0 1 - 0 ---------- --- -    | # rlwinm s2,s2,8,0,31 	-skip_c
| 1001001000    | 01010000001000101100000000001110 0 0 0 - ---  1 1 1 -  0 00 00 00 00 0 0  0 1 - 0 ---------- --- -    | # rlwimi s2,s1,24,0,7 	-skip_c
| 1001001010    | 001110-------------------------- 1 - 0 - ---  0 0 - -  0 10 01 01 01 1 1  0 0 - 0 ---------- --- -    | # addi RA,RA,D

| 1001010000    | 011111-----00000-----00000111000 0 0 0 - ---  1 0 0 -  0 11 00 01 00 0 0  0 0 - 0 ---------- --- -    | # and s0,RB,RB 	-lfsx,lfsux
| 1001010010    | 00111000000000000000000000000001 0 0 1 0 111  1 1 - -  0 00 00 00 00 0 0  0 0 0 0 ---------- 010 -    | # addi s0,s0,1 	-loop_begin,cnt=3
| 1001010100    | 01111100001-----000000001010111- 0 0 0 0 ---  1 0 1 -  0 00 01 00 00 0 -  0 0 - 0 ---------- --- -    | # lbzx s1,RA,s0
| 1001010110    | 01010100010000100100000000111110 0 0 0 - ---  1 1 - -  0 00 00 00 00 0 0  0 1 - 0 ---------- --- -    | # rlwinm s2,s2,8,0,31 	-skip_c
| 1001011000    | 01010000001000101100000000001110 0 0 0 - ---  1 1 1 -  0 00 00 00 00 0 0  0 1 - 0 ---------- --- -    | # rlwimi s2,s1,24,0,7 	-skip_c
| 1001011010    | 00111000001-----1111111111111101 0 - 0 - ---  1 0 - -  0 00 01 00 00 0 0  0 0 - 0 ---------- --- -    | # addi s1,RA,-3

| 1010000000    | 00111000000--------------------- 0 0 0 - ---  1 0 - -  0 00 01 01 01 1 1  0 0 - 0 ---------- --- -    | # addi s0,RA,D 	-lfd,lfdu
| 1010000010    | 00111000000000000000000000000001 0 0 1 0 111  1 1 - -  0 00 00 00 00 0 0  0 0 0 0 ---------- 110 -    | # addi s0,s0,1 	-loop_begin,cnt=7
| 1010000100    | 10001000001000000000000000000000 0 0 0 0 ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # lbz s1,0(s0)
| 1010000110    | 01111000010000101100000000000010 0 0 1 0 111  1 1 - -  0 00 00 00 00 0 0  0 1 0 0 ---------- 110 -    | # rldicl s2,s2,56,0 	-skip_c,loop_begin,cnt=7
| 1010001000    | 01010000010000010000011000111110 0 0 0 1 ---  1 1 1 -  0 00 00 00 00 0 0  0 1 - 0 ---------- --- -    | # rlwimi s1,s2,0,24,31 	-skip_c,loop_end
| 1010001010    | 01111100000000000001010011111110 0 1 0 - ---  0 - 1 -  0 01 00 00 00 0 0  0 0 - 0 ---------- --- -    | # mffgpr RT,s2,0 	-end for non-update

| 1010010000    | 011111-----00000-----00000111000 0 0 0 - ---  1 0 0 -  0 11 00 01 00 0 0  0 0 - 0 ---------- --- 0    | # and s0,RB,RB 	-lfdx,lfdux,lfdepx
| 1010010010    | 00111000000000000000000000000001 0 0 1 0 111  1 1 - -  0 00 00 00 00 0 0  0 0 0 0 ---------- 110 0    | # addi s0,s0,1 	-loop_begin,cnt=7
| 1010010100    | 01111100001-----000000001010111- 0 0 0 0 ---  1 0 1 -  0 00 01 00 00 0 -  0 0 - 0 ---------- --- 1    | # lbzx s1,RA,s0
| 1010010110    | 01111000010000101100000000000010 0 0 1 0 111  1 1 - -  0 00 00 00 00 0 0  0 1 0 0 ---------- 110 0    | # rldicl s2,s2,56,0 	-skip_c,loop_begin,cnt=7
| 1010011000    | 01010000010000010000011000111110 0 0 0 1 ---  1 1 1 -  0 00 00 00 00 0 0  0 1 - 0 ---------- --- 0    | # rlwimi s1,s2,0,24,31 	-skip_c,loop_end
| 1010011010    | 011111-----000000001010011111110 0 1 0 - ---  0 - 1 -  0 01 00 00 00 0 0  0 0 - 0 ---------- --- 0    | # mffgpr RT,s2,0 	-end for non-update
| 1010011100    | 011111-----000010000001000010100 1 - 0 - ---  0 1 1 -  0 10 00 00 00 0 0  0 0 - 0 ---------- --- 0    | # add RA,s1,s0

| 1100110000    | 0111110000100000-----10110111010 0 - 0 - ---  1 - 0 -  0 00 00 10 00 0 0  0 0 - 0 ---------- --- -    | # mfitgpr s1,FRS 	-stfiwx
| 1100110010    | 01010100001000100100000000111110 0 - 0 - ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # rlwinm s2,s1,8,0,31
| 1100110100    | 01010000010000101000010000101110 0 - 0 - ---  1 1 1 -  0 00 00 00 00 0 0  0 1 - 0 ---------- --- -    | # rlwimi s2,s2,16,16,23 	-skip_c
| 1100110110    | 0111110001000000-----0011010111- 0 - 1 0 111  - 1 0 1  0 00 00 01 00 0 -  0 0 0 0 ---------- 010 -    | # stbx s2,s0,RB 	-loop_begin,cnt=3
| 1100111000    | 01010100010000100100000000111110 0 - 0 1 ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # rlwinm s2,s2,8,0,31 	-loop_end

| 1101000000    | 0111110000100000-----10111111100 0 0 0 - ---  1 - 0 -  0 00 00 10 00 0 0  0 0 - 0 ---------- --- -    | # mfstgpr s1,FRS	-stfs,stfsu
| 1101000010    | 01010100001000100100000000111110 0 0 0 - ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # rlwinm s2,s1,8,0,31
| 1101000100    | 01010000010000101000010000101110 0 0 0 - ---  1 1 1 -  0 00 00 00 00 0 0  0 1 - 0 ---------- --- -    | # rlwimi s2,s2,16,16,23 	-skip_c
| 1101000110    | 10011000010000000000000000000000 0 0 1 0 111  - 1 - 1  0 00 00 00 00 0 0  0 0 0 0 ---------- 010 -    | # stb s2,0(s0) 	-loop_begin,cnt=3
| 1101001000    | 01010100010000100100000000111110 0 0 0 1 ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # rlwinm s2,s2,8,0,31 	-loop_end
| 1101001010    | 001110-------------------------- 1 - 0 - ---  0 0 - -  0 10 01 01 01 1 1  0 0 - 0 ---------- --- -    | # addi RA,RA,D

| 1101010000    | 0111110000100000-----10111111100 0 0 0 - ---  1 - 0 -  0 00 00 10 00 0 0  0 0 - 0 ---------- --- -    | # mfstgpr s1,FRS	-stfsx,stfsux
| 1101010010    | 01010100001000100100000000111110 0 0 0 - ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # rlwinm s2,s1,8,0,31
| 1101010100    | 01010000010000101000010000101110 0 0 0 - ---  1 1 1 -  0 00 00 00 00 0 0  0 1 - 0 ---------- --- -    | # rlwimi s2,s2,16,16,23 	-skip_c
| 1101010110    | 0111110001000000-----0011010111- 0 0 1 0 111  - 1 0 1  0 00 00 01 00 0 -  0 0 0 0 ---------- 010 -    | # stbx s2,s0,RB 	-loop_begin,cnt=3
| 1101011000    | 01010100010000100100000000111110 0 0 0 1 ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # rlwinm s2,s2,8,0,31 	-loop_end
| 1101011010    | 011111---------------01000010100 1 - 0 - ---  0 0 0 -  0 10 01 01 00 0 0  0 0 - 0 ---------- --- -    | # add RA,RA,RB

| 1110000000    | 0111110000100000-----10111111110 0 0 0 - ---  1 - 0 -  0 00 00 10 00 0 0  0 0 - 0 ---------- --- -    | # mftgpr s1,FRS 	-stfd,stfdu
| 1110000010    | 01111000010000101100000000000010 0 0 1 0 111  1 1 - -  0 00 00 00 00 0 0  0 1 0 0 ---------- 111 -    | # rldicl s2,s2,56,0 	-skip_c,loop_begin,cnt=8
| 1110000100    | 01010000010000010000011000111110 0 0 0 1 ---  1 1 1 -  0 00 00 00 00 0 0  0 1 - 0 ---------- --- -    | # rlwimi s1,s2,0,24,31 	-skip_c,loop_end
| 1110000110    | 00111000000-----0000000000000000 0 0 0 - ---  1 0 - -  0 00 01 00 00 0 0  0 0 - 0 ---------- --- -    | # addi s0,RA,0
| 1110001000    | 00111000000000000000000000000001 0 0 1 0 111  1 1 - -  0 00 00 00 00 0 0  0 0 0 0 ---------- 110 -    | # addi s0,s0,1 	-loop_begin,cnt=7
| 1110001010    | 1001100001000000---------------- 0 1 0 1 ---  - 1 - 1  0 00 00 01 01 1 1  0 0 - 0 ---------- --- -    | # stb s2,D(s0) 	-loop_end,end for non-update

| 1110010000    | 0111110000100000-----10111111110 0 0 0 - ---  1 - 0 -  0 00 00 10 00 0 0  0 0 - 0 ---------- --- 0    | # mftgpr s1,FRS 	-stfdx,stfdux,stfdepx
| 1110010010    | 01111000010000101100000000000010 0 0 1 0 111  1 1 - -  0 00 00 00 00 0 0  0 1 0 0 ---------- 111 0    | # rldicl s2,s2,56,0 	-skip_c,loop_begin,cnt=8
| 1110010100    | 01010000010000010000011000111110 0 0 0 1 ---  1 1 1 -  0 00 00 00 00 0 0  0 1 - 0 ---------- --- 0    | # rlwimi s1,s2,0,24,31 	-skip_c,loop_end
| 1110010110    | 00111000000-----0000000000000000 0 0 0 - ---  1 0 - -  0 00 01 00 00 0 0  0 0 - 0 ---------- --- 0    | # addi s0,RA,0
| 1110011000    | 00111000000000000000000000000001 0 0 1 0 111  1 1 - -  0 00 00 00 00 0 0  0 0 0 0 ---------- 110 0    | # addi s0,s0,1 	-loop_begin,cnt=7
| 1110011010    | 0111110001000000-----0011010111- 0 1 0 1 ---  - 1 0 1  0 00 00 01 00 0 -  0 0 - 0 ---------- --- 1    | # stbx s2,s0,RB 	-loop_end,end for non-update



| 1111000000    | 110000-------------------------- 0 - 0 - ---  0 0 - -  0 01 01 01 01 1 1  0 0 - 0 ---------- --- -    | # lfs FRT,DS(RA) 	-lfsu

| 1111001000    | 01111100000----------01000010100 0 - 0 - ---  1 0 0 -  0 00 01 01 00 0 0  0 0 - 0 ---------- --- -    | # add s0,RA,RB 	-lfsux
| 1111001010    | 01101000000-----0000000000000000 1 - 0 - ---  0 1 - -  0 00 01 00 00 0 0  0 0 - 0 ---------- --- -    | # xori RA,s0,0

| 1111010000    | 110010-------------------------- 0 - 0 - ---  0 0 - -  0 01 01 01 01 1 1  0 0 - 0 ---------- --- -    | # lfd FRT,DS(RA) 	-lfdu

| 1111011000    | 01111100000----------01000010100 0 - 0 - ---  1 0 0 -  0 00 01 01 00 0 0  0 0 - 0 ---------- --- -    | # add s0,RA,RB 	-lfdux
| 1111011010    | 01101000000-----0000000000000000 1 - 0 - ---  0 1 - -  0 00 01 00 00 0 0  0 0 - 0 ---------- --- -    | # xori RA,s0,0


| 1100000000    | 11111100001---------------100000 0 - 0 - ---  1 - 0 -  0 00 -- 01 -- 0 0  0 0 - 0 ---------- --- -    | # prenrm s1,FB         - prenorm both DP, SP

| 1100001000    | 11111100001---------------100000 0 - 0 - ---  1 - 0 -  0 00 -- 01 -- 0 0  0 0 - 0 ---------- --- -    | # prenrm s1,FB         - prenorm both DP, SP
| 1100001010    | -----------0001000001----------- 1 - 0 - ---  0 1 1 0  1 01 00 00 01 1 1  0 0 - 0 ---------- --- -    | # vvvvv FT,s2,FC,s1    - Original qpx op except B

| 1100010000    | 11101100001---------------100000 0 - 0 - ---  1 - 0 -  0 00 -- 01 -- 0 0  0 0 - 0 ---------- --- -    | # prenrm s1,FB         - prenorm SP only
*END*===========+=======================================================================================================+
?TABLE END rom_instr;
*/


assign rom_instr_pt[1] =
    (({ rom_addr_l2[1] , rom_addr_l2[3] , 
    rom_addr_l2[4] , rom_addr_l2[5] , 
    rom_addr_l2[6] , rom_addr_l2[7] , 
    rom_addr_l2[8] }) === 7'b0000000);
assign rom_instr_pt[2] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] , 
    rom_addr_l2[4] , rom_addr_l2[5] , 
    rom_addr_l2[6] , rom_addr_l2[7] , 
    rom_addr_l2[8] }) === 7'b0000000);
assign rom_instr_pt[3] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] , 
    rom_addr_l2[4] , rom_addr_l2[5] , 
    rom_addr_l2[6] , rom_addr_l2[7] , 
    rom_addr_l2[8] }) === 7'b1010000);
assign rom_instr_pt[4] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] , 
    rom_addr_l2[5] , rom_addr_l2[6] , 
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 6'b000000);
assign rom_instr_pt[5] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] , 
    rom_addr_l2[5] , rom_addr_l2[6] , 
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 6'b100000);
assign rom_instr_pt[6] =
    (({ rom_addr_l2[1] , rom_addr_l2[3] , 
    rom_addr_l2[4] , rom_addr_l2[5] , 
    rom_addr_l2[6] , rom_addr_l2[7] , 
    rom_addr_l2[8] }) === 7'b0001000);
assign rom_instr_pt[7] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] , 
    rom_addr_l2[3] , rom_addr_l2[4] , 
    rom_addr_l2[5] , rom_addr_l2[6] , 
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 8'b11101000);
assign rom_instr_pt[8] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] , 
    rom_addr_l2[3] , rom_addr_l2[4] , 
    rom_addr_l2[5] , rom_addr_l2[6] , 
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 8'b10111000);
assign rom_instr_pt[9] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] , 
    rom_addr_l2[3] , rom_addr_l2[5] , 
    rom_addr_l2[6] , rom_addr_l2[7] , 
    rom_addr_l2[8] }) === 7'b0011000);
assign rom_instr_pt[10] =
    (({ rom_addr_l2[0] , rom_addr_l2[2] , 
    rom_addr_l2[5] , rom_addr_l2[6] , 
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 6'b011000);
assign rom_instr_pt[11] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] , 
    rom_addr_l2[3] , rom_addr_l2[4] , 
    rom_addr_l2[6] , rom_addr_l2[7] , 
    rom_addr_l2[8] }) === 7'b0100000);
assign rom_instr_pt[12] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] , 
    rom_addr_l2[2] , rom_addr_l2[4] , 
    rom_addr_l2[6] , rom_addr_l2[7] , 
    rom_addr_l2[8] }) === 7'b0100000);
assign rom_instr_pt[13] =
    (({ rom_addr_l2[0] , rom_addr_l2[3] , 
    rom_addr_l2[4] , rom_addr_l2[6] , 
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 6'b001000);
assign rom_instr_pt[14] =
    (({ rom_addr_l2[2] , rom_addr_l2[3] , 
    rom_addr_l2[4] , rom_addr_l2[6] , 
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 6'b111000);
assign rom_instr_pt[15] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] , 
    rom_addr_l2[4] , rom_addr_l2[6] , 
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 6'b101000);
assign rom_instr_pt[16] =
    (({ rom_addr_l2[0] , rom_addr_l2[2] , 
    rom_addr_l2[4] , rom_addr_l2[6] , 
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 6'b101000);
assign rom_instr_pt[17] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] , 
    rom_addr_l2[4] , rom_addr_l2[6] , 
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 6'b111000);
assign rom_instr_pt[18] =
    (({ rom_addr_l2[0] , rom_addr_l2[4] , 
    rom_addr_l2[6] , rom_addr_l2[7] , 
    rom_addr_l2[8] }) === 5'b01000);
assign rom_instr_pt[19] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] , 
    rom_addr_l2[2] , rom_addr_l2[3] , 
    rom_addr_l2[6] , rom_addr_l2[7] , 
    rom_addr_l2[8] }) === 7'b1000000);
assign rom_instr_pt[20] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] , 
    rom_addr_l2[2] , rom_addr_l2[3] , 
    rom_addr_l2[6] , rom_addr_l2[7] , 
    rom_addr_l2[8] }) === 7'b1110000);
assign rom_instr_pt[21] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] , 
    rom_addr_l2[2] , rom_addr_l2[3] , 
    rom_addr_l2[6] , rom_addr_l2[7] , 
    rom_addr_l2[8] }) === 7'b1101000);
assign rom_instr_pt[22] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] , 
    rom_addr_l2[6] , rom_addr_l2[7] , 
    rom_addr_l2[8] }) === 5'b11000);
assign rom_instr_pt[23] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] , 
    rom_addr_l2[3] , rom_addr_l2[4] , 
    rom_addr_l2[6] , rom_addr_l2[7] , 
    rom_addr_l2[8] }) === 7'b0100100);
assign rom_instr_pt[24] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] , 
    rom_addr_l2[2] , rom_addr_l2[4] , 
    rom_addr_l2[6] , rom_addr_l2[7] , 
    rom_addr_l2[8] }) === 7'b0011100);
assign rom_instr_pt[25] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] , 
    rom_addr_l2[2] , rom_addr_l2[3] , 
    rom_addr_l2[6] , rom_addr_l2[7] , 
    rom_addr_l2[8] }) === 7'b0011100);
assign rom_instr_pt[26] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] , 
    rom_addr_l2[3] , rom_addr_l2[6] , 
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 6'b011100);
assign rom_instr_pt[27] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] , 
    rom_addr_l2[2] , rom_addr_l2[3] , 
    rom_addr_l2[6] , rom_addr_l2[7] , 
    rom_addr_l2[8] }) === 7'b0111100);
assign rom_instr_pt[28] =
    (({ rom_addr_l2[0] , rom_addr_l2[2] , 
    rom_addr_l2[6] , rom_addr_l2[7] , 
    rom_addr_l2[8] }) === 5'b01100);
assign rom_instr_pt[29] =
    (({ rom_addr_l2[0] , rom_addr_l2[3] , 
    rom_addr_l2[4] , rom_addr_l2[5] , 
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 6'b001000);
assign rom_instr_pt[30] =
    (({ rom_addr_l2[0] , rom_addr_l2[2] , 
    rom_addr_l2[3] , rom_addr_l2[4] , 
    rom_addr_l2[5] , rom_addr_l2[7] , 
    rom_addr_l2[8] }) === 7'b0111100);
assign rom_instr_pt[31] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] , 
    rom_addr_l2[2] , rom_addr_l2[3] , 
    rom_addr_l2[4] , rom_addr_l2[7] , 
    rom_addr_l2[8] }) === 7'b0110000);
assign rom_instr_pt[32] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] , 
    rom_addr_l2[3] , rom_addr_l2[4] , 
    rom_addr_l2[5] , rom_addr_l2[6] , 
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 8'b01001010);
assign rom_instr_pt[33] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] , 
    rom_addr_l2[4] , rom_addr_l2[5] , 
    rom_addr_l2[6] , rom_addr_l2[7] , 
    rom_addr_l2[8] }) === 7'b0111010);
assign rom_instr_pt[34] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] , 
    rom_addr_l2[3] , rom_addr_l2[4] , 
    rom_addr_l2[6] , rom_addr_l2[7] , 
    rom_addr_l2[8] }) === 7'b0110010);
assign rom_instr_pt[35] =
    (({ rom_addr_l2[1] , rom_addr_l2[4] , 
    rom_addr_l2[6] , rom_addr_l2[7] , 
    rom_addr_l2[8] }) === 5'b10110);
assign rom_instr_pt[36] =
    (({ rom_addr_l2[1] , rom_addr_l2[4] , 
    rom_addr_l2[6] , rom_addr_l2[7] , 
    rom_addr_l2[8] }) === 5'b01110);
assign rom_instr_pt[37] =
    (({ rom_addr_l2[1] , rom_addr_l2[3] , 
    rom_addr_l2[6] , rom_addr_l2[7] , 
    rom_addr_l2[8] }) === 5'b10110);
assign rom_instr_pt[38] =
    (({ rom_addr_l2[2] , rom_addr_l2[3] , 
    rom_addr_l2[6] , rom_addr_l2[7] , 
    rom_addr_l2[8] }) === 5'b11110);
assign rom_instr_pt[39] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] , 
    rom_addr_l2[3] , rom_addr_l2[4] , 
    rom_addr_l2[5] , rom_addr_l2[7] , 
    rom_addr_l2[8] }) === 7'b0110010);
assign rom_instr_pt[40] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] , 
    rom_addr_l2[4] , rom_addr_l2[5] , 
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 6'b010010);
assign rom_instr_pt[41] =
    (({ rom_addr_l2[1] , rom_addr_l2[4] , 
    rom_addr_l2[5] , rom_addr_l2[7] , 
    rom_addr_l2[8] }) === 5'b00010);
assign rom_instr_pt[42] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] , 
    rom_addr_l2[3] , rom_addr_l2[4] , 
    rom_addr_l2[5] , rom_addr_l2[7] , 
    rom_addr_l2[8] }) === 7'b0011010);
assign rom_instr_pt[43] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] , 
    rom_addr_l2[3] , rom_addr_l2[5] , 
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 6'b000010);
assign rom_instr_pt[44] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] , 
    rom_addr_l2[3] , rom_addr_l2[5] , 
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 6'b001010);
assign rom_instr_pt[45] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] , 
    rom_addr_l2[2] , rom_addr_l2[3] , 
    rom_addr_l2[5] , rom_addr_l2[7] , 
    rom_addr_l2[8] }) === 7'b0000110);
assign rom_instr_pt[46] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] , 
    rom_addr_l2[2] , rom_addr_l2[3] , 
    rom_addr_l2[5] , rom_addr_l2[7] , 
    rom_addr_l2[8] }) === 7'b0100110);
assign rom_instr_pt[47] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] , 
    rom_addr_l2[3] , rom_addr_l2[5] , 
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 6'b001110);
assign rom_instr_pt[48] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] , 
    rom_addr_l2[3] , rom_addr_l2[4] , 
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 6'b110010);
assign rom_instr_pt[49] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] , 
    rom_addr_l2[2] , rom_addr_l2[3] , 
    rom_addr_l2[4] , rom_addr_l2[7] , 
    rom_addr_l2[8] }) === 7'b0101010);
assign rom_instr_pt[50] =
    (({ rom_addr_l2[2] , rom_addr_l2[3] , 
    rom_addr_l2[4] , rom_addr_l2[7] , 
    rom_addr_l2[8] }) === 5'b11010);
assign rom_instr_pt[51] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] , 
    rom_addr_l2[3] , rom_addr_l2[4] , 
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 6'b111110);
assign rom_instr_pt[52] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] , 
    rom_addr_l2[4] , rom_addr_l2[7] , 
    rom_addr_l2[8] }) === 5'b10110);
assign rom_instr_pt[53] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] , 
    rom_addr_l2[2] , rom_addr_l2[7] , 
    rom_addr_l2[8] }) === 5'b11010);
assign rom_instr_pt[54] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] , 
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 4'b1110);
assign rom_instr_pt[55] =
    (({ rom_addr_l2[1] , rom_addr_l2[3] , 
    rom_addr_l2[4] , rom_addr_l2[6] , 
    rom_addr_l2[8] }) === 5'b10000);
assign rom_instr_pt[56] =
    (({ rom_addr_l2[1] , rom_addr_l2[4] , 
    rom_addr_l2[5] , rom_addr_l2[6] , 
    rom_addr_l2[8] }) === 5'b11010);
assign rom_instr_pt[57] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] , 
    rom_addr_l2[3] , rom_addr_l2[4] , 
    rom_addr_l2[6] , rom_addr_l2[8]
     }) === 6'b100010);
assign rom_instr_pt[58] =
    (({ rom_addr_l2[2] , rom_addr_l2[3] , 
    rom_addr_l2[4] , rom_addr_l2[6] , 
    rom_addr_l2[8] }) === 5'b01010);
assign rom_instr_pt[59] =
    (({ rom_addr_l2[1] , rom_addr_l2[3] , 
    rom_addr_l2[4] , rom_addr_l2[6] , 
    rom_addr_l2[8] }) === 5'b10110);
assign rom_instr_pt[60] =
    (({ rom_addr_l2[1] , rom_addr_l2[3] , 
    rom_addr_l2[4] , rom_addr_l2[6] , 
    rom_addr_l2[8] }) === 5'b11110);
assign rom_instr_pt[61] =
    (({ rom_addr_l2[0] , rom_addr_l2[2] , 
    rom_addr_l2[4] , rom_addr_l2[6] , 
    rom_addr_l2[8] }) === 5'b11110);
assign rom_instr_pt[62] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] , 
    rom_addr_l2[2] , rom_addr_l2[3] , 
    rom_addr_l2[6] , rom_addr_l2[8]
     }) === 6'b111010);
assign rom_instr_pt[63] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] , 
    rom_addr_l2[3] , rom_addr_l2[6] , 
    rom_addr_l2[8] }) === 5'b00110);
assign rom_instr_pt[64] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] , 
    rom_addr_l2[2] , rom_addr_l2[3] , 
    rom_addr_l2[6] , rom_addr_l2[8]
     }) === 6'b110110);
assign rom_instr_pt[65] =
    (({ rom_addr_l2[0] , rom_addr_l2[2] , 
    rom_addr_l2[3] , rom_addr_l2[6] , 
    rom_addr_l2[8] }) === 5'b11110);
assign rom_instr_pt[66] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] , 
    rom_addr_l2[2] , rom_addr_l2[3] , 
    rom_addr_l2[4] , rom_addr_l2[5] , 
    rom_addr_l2[8] }) === 7'b0011000);
assign rom_instr_pt[67] =
    (({ rom_addr_l2[0] , rom_addr_l2[2] , 
    rom_addr_l2[3] , rom_addr_l2[4] , 
    rom_addr_l2[5] , rom_addr_l2[8]
     }) === 6'b011000);
assign rom_instr_pt[68] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] , 
    rom_addr_l2[3] , rom_addr_l2[4] , 
    rom_addr_l2[5] , rom_addr_l2[8]
     }) === 6'b111100);
assign rom_instr_pt[69] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] , 
    rom_addr_l2[3] , rom_addr_l2[8]
     }) === 4'b1100);
assign rom_instr_pt[70] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] , 
    rom_addr_l2[4] , rom_addr_l2[5] , 
    rom_addr_l2[6] , rom_addr_l2[7] , 
    rom_addr_l2[8] }) === 7'b1010001);
assign rom_instr_pt[71] =
    (({ rom_addr_l2[2] , rom_addr_l2[4] , 
    rom_addr_l2[5] , rom_addr_l2[6] , 
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 6'b101001);
assign rom_instr_pt[72] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] , 
    rom_addr_l2[4] , rom_addr_l2[5] , 
    rom_addr_l2[6] , rom_addr_l2[7] , 
    rom_addr_l2[8] }) === 7'b0111001);
assign rom_instr_pt[73] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] , 
    rom_addr_l2[4] , rom_addr_l2[5] , 
    rom_addr_l2[6] , rom_addr_l2[7] , 
    rom_addr_l2[8] }) === 7'b1111001);
assign rom_instr_pt[74] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] , 
    rom_addr_l2[3] , rom_addr_l2[5] , 
    rom_addr_l2[6] , rom_addr_l2[7] , 
    rom_addr_l2[8] }) === 7'b0111001);
assign rom_instr_pt[75] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] , 
    rom_addr_l2[3] , rom_addr_l2[4] , 
    rom_addr_l2[6] , rom_addr_l2[7] , 
    rom_addr_l2[8] }) === 7'b1100001);
assign rom_instr_pt[76] =
    (({ rom_addr_l2[2] , rom_addr_l2[3] , 
    rom_addr_l2[4] , rom_addr_l2[6] , 
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 6'b100001);
assign rom_instr_pt[77] =
    (({ rom_addr_l2[1] , rom_addr_l2[3] , 
    rom_addr_l2[4] , rom_addr_l2[6] , 
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 6'b000001);
assign rom_instr_pt[78] =
    (({ rom_addr_l2[1] , rom_addr_l2[3] , 
    rom_addr_l2[4] , rom_addr_l2[6] , 
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 6'b100001);
assign rom_instr_pt[79] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] , 
    rom_addr_l2[3] , rom_addr_l2[4] , 
    rom_addr_l2[6] , rom_addr_l2[7] , 
    rom_addr_l2[8] }) === 7'b1110001);
assign rom_instr_pt[80] =
    (({ rom_addr_l2[2] , rom_addr_l2[3] , 
    rom_addr_l2[6] , rom_addr_l2[7] , 
    rom_addr_l2[8] }) === 5'b10001);
assign rom_instr_pt[81] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] , 
    rom_addr_l2[3] , rom_addr_l2[6] , 
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 6'b001001);
assign rom_instr_pt[82] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] , 
    rom_addr_l2[6] , rom_addr_l2[7] , 
    rom_addr_l2[8] }) === 5'b00001);
assign rom_instr_pt[83] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] , 
    rom_addr_l2[2] , rom_addr_l2[6] , 
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 6'b110001);
assign rom_instr_pt[84] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] , 
    rom_addr_l2[2] , rom_addr_l2[4] , 
    rom_addr_l2[6] , rom_addr_l2[7] , 
    rom_addr_l2[8] }) === 7'b0011101);
assign rom_instr_pt[85] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] , 
    rom_addr_l2[3] , rom_addr_l2[6] , 
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 6'b000101);
assign rom_instr_pt[86] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] , 
    rom_addr_l2[3] , rom_addr_l2[6] , 
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 6'b010101);
assign rom_instr_pt[87] =
    (({ rom_addr_l2[3] , rom_addr_l2[6] , 
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 4'b0101);
assign rom_instr_pt[88] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] , 
    rom_addr_l2[2] , rom_addr_l2[3] , 
    rom_addr_l2[6] , rom_addr_l2[7] , 
    rom_addr_l2[8] }) === 7'b0011101);
assign rom_instr_pt[89] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] , 
    rom_addr_l2[2] , rom_addr_l2[3] , 
    rom_addr_l2[6] , rom_addr_l2[7] , 
    rom_addr_l2[8] }) === 7'b0111101);
assign rom_instr_pt[90] =
    (({ rom_addr_l2[2] , rom_addr_l2[3] , 
    rom_addr_l2[6] , rom_addr_l2[7] , 
    rom_addr_l2[8] }) === 5'b11101);
assign rom_instr_pt[91] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] , 
    rom_addr_l2[3] , rom_addr_l2[5] , 
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 6'b000001);
assign rom_instr_pt[92] =
    (({ rom_addr_l2[0] , rom_addr_l2[2] , 
    rom_addr_l2[3] , rom_addr_l2[4] , 
    rom_addr_l2[5] , rom_addr_l2[7] , 
    rom_addr_l2[8] }) === 7'b0001101);
assign rom_instr_pt[93] =
    (({ rom_addr_l2[0] , rom_addr_l2[2] , 
    rom_addr_l2[3] , rom_addr_l2[4] , 
    rom_addr_l2[5] , rom_addr_l2[7] , 
    rom_addr_l2[8] }) === 7'b0111101);
assign rom_instr_pt[94] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] , 
    rom_addr_l2[2] , rom_addr_l2[3] , 
    rom_addr_l2[4] , rom_addr_l2[7] , 
    rom_addr_l2[8] }) === 7'b0101001);
assign rom_instr_pt[95] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] , 
    rom_addr_l2[2] , rom_addr_l2[4] , 
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 6'b010001);
assign rom_instr_pt[96] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] , 
    rom_addr_l2[2] , rom_addr_l2[4] , 
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 6'b100101);
assign rom_instr_pt[97] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] , 
    rom_addr_l2[2] , rom_addr_l2[3] , 
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 6'b010001);
assign rom_instr_pt[98] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] , 
    rom_addr_l2[3] , rom_addr_l2[7] , 
    rom_addr_l2[8] }) === 5'b00101);
assign rom_instr_pt[99] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] , 
    rom_addr_l2[2] , rom_addr_l2[7] , 
    rom_addr_l2[8] }) === 5'b10001);
assign rom_instr_pt[100] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] , 
    rom_addr_l2[2] , rom_addr_l2[4] , 
    rom_addr_l2[5] , rom_addr_l2[6] , 
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 8'b01101011);
assign rom_instr_pt[101] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] , 
    rom_addr_l2[3] , rom_addr_l2[4] , 
    rom_addr_l2[6] , rom_addr_l2[7] , 
    rom_addr_l2[8] }) === 7'b1110011);
assign rom_instr_pt[102] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] , 
    rom_addr_l2[4] , rom_addr_l2[6] , 
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 6'b011011);
assign rom_instr_pt[103] =
    (({ rom_addr_l2[2] , rom_addr_l2[3] , 
    rom_addr_l2[6] , rom_addr_l2[7] , 
    rom_addr_l2[8] }) === 5'b11011);
assign rom_instr_pt[104] =
    (({ rom_addr_l2[1] , rom_addr_l2[4] , 
    rom_addr_l2[6] , rom_addr_l2[7] , 
    rom_addr_l2[8] }) === 5'b10111);
assign rom_instr_pt[105] =
    (({ rom_addr_l2[1] , rom_addr_l2[3] , 
    rom_addr_l2[6] , rom_addr_l2[7] , 
    rom_addr_l2[8] }) === 5'b10111);
assign rom_instr_pt[106] =
    (({ rom_addr_l2[1] , rom_addr_l2[3] , 
    rom_addr_l2[6] , rom_addr_l2[7] , 
    rom_addr_l2[8] }) === 5'b01111);
assign rom_instr_pt[107] =
    (({ rom_addr_l2[2] , rom_addr_l2[6] , 
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 4'b0111);
assign rom_instr_pt[108] =
    (({ rom_addr_l2[1] , rom_addr_l2[6] , 
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 4'b0111);
assign rom_instr_pt[109] =
    (({ rom_addr_l2[3] , rom_addr_l2[4] , 
    rom_addr_l2[5] , rom_addr_l2[7] , 
    rom_addr_l2[8] }) === 5'b01011);
assign rom_instr_pt[110] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] , 
    rom_addr_l2[3] , rom_addr_l2[5] , 
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 6'b000011);
assign rom_instr_pt[111] =
    (({ rom_addr_l2[2] , rom_addr_l2[3] , 
    rom_addr_l2[5] , rom_addr_l2[7] , 
    rom_addr_l2[8] }) === 5'b00011);
assign rom_instr_pt[112] =
    (({ rom_addr_l2[1] , rom_addr_l2[3] , 
    rom_addr_l2[5] , rom_addr_l2[7] , 
    rom_addr_l2[8] }) === 5'b00011);
assign rom_instr_pt[113] =
    (({ rom_addr_l2[1] , rom_addr_l2[3] , 
    rom_addr_l2[5] , rom_addr_l2[7] , 
    rom_addr_l2[8] }) === 5'b01011);
assign rom_instr_pt[114] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] , 
    rom_addr_l2[2] , rom_addr_l2[5] , 
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 6'b110011);
assign rom_instr_pt[115] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] , 
    rom_addr_l2[2] , rom_addr_l2[5] , 
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 6'b011011);
assign rom_instr_pt[116] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] , 
    rom_addr_l2[3] , rom_addr_l2[4] , 
    rom_addr_l2[5] , rom_addr_l2[7] , 
    rom_addr_l2[8] }) === 7'b0100111);
assign rom_instr_pt[117] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] , 
    rom_addr_l2[2] , rom_addr_l2[3] , 
    rom_addr_l2[5] , rom_addr_l2[7] , 
    rom_addr_l2[8] }) === 7'b0000111);
assign rom_instr_pt[118] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] , 
    rom_addr_l2[5] , rom_addr_l2[7] , 
    rom_addr_l2[8] }) === 5'b00111);
assign rom_instr_pt[119] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] , 
    rom_addr_l2[2] , rom_addr_l2[5] , 
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 6'b110111);
assign rom_instr_pt[120] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] , 
    rom_addr_l2[3] , rom_addr_l2[4] , 
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 6'b010011);
assign rom_instr_pt[121] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] , 
    rom_addr_l2[3] , rom_addr_l2[4] , 
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 6'b101011);
assign rom_instr_pt[122] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] , 
    rom_addr_l2[2] , rom_addr_l2[4] , 
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 6'b010011);
assign rom_instr_pt[123] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] , 
    rom_addr_l2[3] , rom_addr_l2[4] , 
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 6'b100111);
assign rom_instr_pt[124] =
    (({ rom_addr_l2[2] , rom_addr_l2[3] , 
    rom_addr_l2[4] , rom_addr_l2[7] , 
    rom_addr_l2[8] }) === 5'b11111);
assign rom_instr_pt[125] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] , 
    rom_addr_l2[3] , rom_addr_l2[7] , 
    rom_addr_l2[8] }) === 5'b10011);
assign rom_instr_pt[126] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] , 
    rom_addr_l2[3] , rom_addr_l2[7] , 
    rom_addr_l2[8] }) === 5'b00111);
assign rom_instr_pt[127] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] , 
    rom_addr_l2[2] , rom_addr_l2[7] , 
    rom_addr_l2[8] }) === 5'b10011);
assign rom_instr_pt[128] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] , 
    rom_addr_l2[2] , rom_addr_l2[7] , 
    rom_addr_l2[8] }) === 5'b11111);
assign rom_instr_pt[129] =
    (({ rom_addr_l2[0] , rom_addr_l2[2] , 
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 4'b1111);
assign rom_instr_pt[130] =
    (({ rom_addr_l2[1] , rom_addr_l2[3] , 
    rom_addr_l2[4] , rom_addr_l2[5] , 
    rom_addr_l2[6] , rom_addr_l2[8]
     }) === 6'b111001);
assign rom_instr_pt[131] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] , 
    rom_addr_l2[3] , rom_addr_l2[4] , 
    rom_addr_l2[5] , rom_addr_l2[6] , 
    rom_addr_l2[8] }) === 7'b0101101);
assign rom_instr_pt[132] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] , 
    rom_addr_l2[3] , rom_addr_l2[4] , 
    rom_addr_l2[6] , rom_addr_l2[8]
     }) === 6'b010001);
assign rom_instr_pt[133] =
    (({ rom_addr_l2[0] , rom_addr_l2[2] , 
    rom_addr_l2[3] , rom_addr_l2[4] , 
    rom_addr_l2[6] , rom_addr_l2[8]
     }) === 6'b010001);
assign rom_instr_pt[134] =
    (({ rom_addr_l2[2] , rom_addr_l2[3] , 
    rom_addr_l2[4] , rom_addr_l2[6] , 
    rom_addr_l2[8] }) === 5'b01001);
assign rom_instr_pt[135] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] , 
    rom_addr_l2[3] , rom_addr_l2[4] , 
    rom_addr_l2[6] , rom_addr_l2[8]
     }) === 6'b011101);
assign rom_instr_pt[136] =
    (({ rom_addr_l2[2] , rom_addr_l2[3] , 
    rom_addr_l2[4] , rom_addr_l2[5] , 
    rom_addr_l2[6] , rom_addr_l2[8]
     }) === 6'b010011);
assign rom_instr_pt[137] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] , 
    rom_addr_l2[3] , rom_addr_l2[5] , 
    rom_addr_l2[6] , rom_addr_l2[8]
     }) === 6'b110011);
assign rom_instr_pt[138] =
    (({ rom_addr_l2[1] , rom_addr_l2[3] , 
    rom_addr_l2[5] , rom_addr_l2[6] , 
    rom_addr_l2[8] }) === 5'b10011);
assign rom_instr_pt[139] =
    (({ rom_addr_l2[2] , rom_addr_l2[5] , 
    rom_addr_l2[6] , rom_addr_l2[8]
     }) === 4'b0011);
assign rom_instr_pt[140] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] , 
    rom_addr_l2[3] , rom_addr_l2[4] , 
    rom_addr_l2[5] , rom_addr_l2[6] , 
    rom_addr_l2[8] }) === 7'b0100111);
assign rom_instr_pt[141] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] , 
    rom_addr_l2[3] , rom_addr_l2[5] , 
    rom_addr_l2[6] , rom_addr_l2[8]
     }) === 6'b110111);
assign rom_instr_pt[142] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] , 
    rom_addr_l2[5] , rom_addr_l2[6] , 
    rom_addr_l2[8] }) === 5'b00111);
assign rom_instr_pt[143] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] , 
    rom_addr_l2[2] , rom_addr_l2[5] , 
    rom_addr_l2[6] , rom_addr_l2[8]
     }) === 6'b110111);
assign rom_instr_pt[144] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] , 
    rom_addr_l2[3] , rom_addr_l2[4] , 
    rom_addr_l2[6] , rom_addr_l2[8]
     }) === 6'b000011);
assign rom_instr_pt[145] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] , 
    rom_addr_l2[3] , rom_addr_l2[4] , 
    rom_addr_l2[6] , rom_addr_l2[8]
     }) === 6'b100011);
assign rom_instr_pt[146] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] , 
    rom_addr_l2[3] , rom_addr_l2[4] , 
    rom_addr_l2[6] , rom_addr_l2[8]
     }) === 6'b010011);
assign rom_instr_pt[147] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] , 
    rom_addr_l2[4] , rom_addr_l2[6] , 
    rom_addr_l2[8] }) === 5'b11111);
assign rom_instr_pt[148] =
    (({ rom_addr_l2[2] , rom_addr_l2[3] , 
    rom_addr_l2[6] , rom_addr_l2[8]
     }) === 4'b0011);
assign rom_instr_pt[149] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] , 
    rom_addr_l2[2] , rom_addr_l2[3] , 
    rom_addr_l2[6] , rom_addr_l2[8]
     }) === 6'b111011);
assign rom_instr_pt[150] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] , 
    rom_addr_l2[2] , rom_addr_l2[3] , 
    rom_addr_l2[6] , rom_addr_l2[8]
     }) === 6'b110111);
assign rom_instr_pt[151] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] , 
    rom_addr_l2[6] , rom_addr_l2[8]
     }) === 4'b0011);
assign rom_instr_pt[152] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] , 
    rom_addr_l2[2] , rom_addr_l2[6] , 
    rom_addr_l2[8] }) === 5'b11011);
assign rom_instr_pt[153] =
    (({ rom_addr_l2[0] , rom_addr_l2[2] , 
    rom_addr_l2[3] , rom_addr_l2[4] , 
    rom_addr_l2[5] , rom_addr_l2[8]
     }) === 6'b011001);
assign rom_instr_pt[154] =
    (({ rom_addr_l2[2] , rom_addr_l2[3] , 
    rom_addr_l2[4] , rom_addr_l2[5] , 
    rom_addr_l2[8] }) === 5'b11001);
assign rom_instr_pt[155] =
    (({ rom_addr_l2[0] , rom_addr_l2[2] , 
    rom_addr_l2[3] , rom_addr_l2[4] , 
    rom_addr_l2[5] , rom_addr_l2[8]
     }) === 6'b010101);
assign rom_instr_pt[156] =
    (({ rom_addr_l2[0] , rom_addr_l2[2] , 
    rom_addr_l2[3] , rom_addr_l2[4] , 
    rom_addr_l2[5] , rom_addr_l2[8]
     }) === 6'b011101);
assign rom_instr_pt[157] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] , 
    rom_addr_l2[2] , rom_addr_l2[4] , 
    rom_addr_l2[5] , rom_addr_l2[8]
     }) === 6'b010111);
assign rom_instr_pt[158] =
    (({ rom_addr_l2[1] , rom_addr_l2[3] , 
    rom_addr_l2[4] , rom_addr_l2[8]
     }) === 4'b1111);
assign rom_instr_pt[159] =
    (({ rom_addr_l2[0] , rom_addr_l2[2] , 
    rom_addr_l2[4] , rom_addr_l2[8]
     }) === 4'b1111);
assign rom_instr_pt[160] =
    (({ rom_addr_l2[0] , rom_addr_l2[2] , 
    rom_addr_l2[3] , rom_addr_l2[8]
     }) === 4'b1111);
assign rom_instr_pt[161] =
    (({ rom_addr_l2[3] , rom_addr_l2[8]
     }) === 2'b11);
assign rom_instr_pt[162] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] , 
    rom_addr_l2[8] }) === 3'b011);
assign rom_instr_pt[163] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] , 
    rom_addr_l2[3] , rom_addr_l2[5] , 
    rom_addr_l2[6] , rom_addr_l2[7]
     }) === 6'b011100);
assign rom_instr_pt[164] =
    (({ rom_addr_l2[2] , rom_addr_l2[3] , 
    rom_addr_l2[4] , rom_addr_l2[6] , 
    rom_addr_l2[7] }) === 5'b10000);
assign rom_instr_pt[165] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] , 
    rom_addr_l2[2] , rom_addr_l2[3] , 
    rom_addr_l2[6] , rom_addr_l2[7]
     }) === 6'b010000);
assign rom_instr_pt[166] =
    (({ rom_addr_l2[0] , rom_addr_l2[2] , 
    rom_addr_l2[3] , rom_addr_l2[4] , 
    rom_addr_l2[5] , rom_addr_l2[7]
     }) === 6'b011100);
assign rom_instr_pt[167] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] , 
    rom_addr_l2[3] , rom_addr_l2[4] , 
    rom_addr_l2[5] , rom_addr_l2[7]
     }) === 6'b000010);
assign rom_instr_pt[168] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] , 
    rom_addr_l2[3] , rom_addr_l2[4] , 
    rom_addr_l2[5] , rom_addr_l2[6] , 
    rom_addr_l2[7] }) === 7'b0101101);
assign rom_instr_pt[169] =
    (({ rom_addr_l2[0] , rom_addr_l2[3] , 
    rom_addr_l2[4] , rom_addr_l2[6] , 
    rom_addr_l2[7] }) === 5'b00101);
assign rom_instr_pt[170] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] , 
    rom_addr_l2[3] , rom_addr_l2[6] , 
    rom_addr_l2[7] }) === 5'b11101);
assign rom_instr_pt[171] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] , 
    rom_addr_l2[3] , rom_addr_l2[6] , 
    rom_addr_l2[7] }) === 5'b01101);
assign rom_instr_pt[172] =
    (({ rom_addr_l2[3] , rom_addr_l2[4] , 
    rom_addr_l2[6] , rom_addr_l2[7]
     }) === 4'b0011);
assign rom_instr_pt[173] =
    (({ rom_addr_l2[1] , rom_addr_l2[4] , 
    rom_addr_l2[6] , rom_addr_l2[7]
     }) === 4'b0111);
assign rom_instr_pt[174] =
    (({ rom_addr_l2[2] , rom_addr_l2[3] , 
    rom_addr_l2[4] , rom_addr_l2[5] , 
    rom_addr_l2[7] }) === 5'b10101);
assign rom_instr_pt[175] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] , 
    rom_addr_l2[4] , rom_addr_l2[5] , 
    rom_addr_l2[7] }) === 5'b10101);
assign rom_instr_pt[176] =
    (({ rom_addr_l2[2] , rom_addr_l2[4] , 
    rom_addr_l2[5] , rom_addr_l2[7]
     }) === 4'b1101);
assign rom_instr_pt[177] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] , 
    rom_addr_l2[3] , rom_addr_l2[5] , 
    rom_addr_l2[7] }) === 5'b10001);
assign rom_instr_pt[178] =
    (({ rom_addr_l2[2] , rom_addr_l2[3] , 
    rom_addr_l2[5] , rom_addr_l2[7]
     }) === 4'b0001);
assign rom_instr_pt[179] =
    (({ rom_addr_l2[2] , rom_addr_l2[3] , 
    rom_addr_l2[5] , rom_addr_l2[7]
     }) === 4'b1101);
assign rom_instr_pt[180] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] , 
    rom_addr_l2[2] , rom_addr_l2[4] , 
    rom_addr_l2[5] , rom_addr_l2[7]
     }) === 6'b010111);
assign rom_instr_pt[181] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] , 
    rom_addr_l2[2] , rom_addr_l2[3] , 
    rom_addr_l2[5] , rom_addr_l2[7]
     }) === 6'b000011);
assign rom_instr_pt[182] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] , 
    rom_addr_l2[2] , rom_addr_l2[3] , 
    rom_addr_l2[5] , rom_addr_l2[7]
     }) === 6'b010011);
assign rom_instr_pt[183] =
    (({ rom_addr_l2[2] , rom_addr_l2[3] , 
    rom_addr_l2[4] , rom_addr_l2[7]
     }) === 4'b1111);
assign rom_instr_pt[184] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] , 
    rom_addr_l2[2] , rom_addr_l2[4] , 
    rom_addr_l2[7] }) === 5'b01011);
assign rom_instr_pt[185] =
    (({ rom_addr_l2[0] , rom_addr_l2[4] , 
    rom_addr_l2[5] , rom_addr_l2[6]
     }) === 4'b1100);
assign rom_instr_pt[186] =
    (({ rom_addr_l2[0] , rom_addr_l2[2] , 
    rom_addr_l2[4] , rom_addr_l2[5] , 
    rom_addr_l2[6] }) === 5'b01110);
assign rom_instr_pt[187] =
    (({ rom_addr_l2[0] , rom_addr_l2[2] , 
    rom_addr_l2[4] , rom_addr_l2[5] , 
    rom_addr_l2[6] }) === 5'b11110);
assign rom_instr_pt[188] =
    (({ rom_addr_l2[3] , rom_addr_l2[5] , 
    rom_addr_l2[6] }) === 3'b010);
assign rom_instr_pt[189] =
    (({ rom_addr_l2[5] , rom_addr_l2[6]
     }) === 2'b10);
assign rom_instr_pt[190] =
    (({ rom_addr_l2[0] , rom_addr_l2[2] , 
    rom_addr_l2[3] , rom_addr_l2[4] , 
    rom_addr_l2[6] }) === 5'b10000);
assign rom_instr_pt[191] =
    (({ rom_addr_l2[0] , rom_addr_l2[2] , 
    rom_addr_l2[4] , rom_addr_l2[6]
     }) === 4'b1110);
assign rom_instr_pt[192] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] , 
    rom_addr_l2[2] , rom_addr_l2[3] , 
    rom_addr_l2[6] }) === 5'b11110);
assign rom_instr_pt[193] =
    (({ rom_addr_l2[0] , rom_addr_l2[2] , 
    rom_addr_l2[3] , rom_addr_l2[6]
     }) === 4'b1110);
assign rom_instr_pt[194] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] , 
    rom_addr_l2[2] , rom_addr_l2[4] , 
    rom_addr_l2[5] , rom_addr_l2[6]
     }) === 6'b010001);
assign rom_instr_pt[195] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] , 
    rom_addr_l2[2] , rom_addr_l2[3] , 
    rom_addr_l2[4] , rom_addr_l2[5] , 
    rom_addr_l2[6] }) === 7'b0101011);
assign rom_instr_pt[196] =
    (({ rom_addr_l2[1] , rom_addr_l2[3] , 
    rom_addr_l2[4] , rom_addr_l2[5] , 
    rom_addr_l2[6] }) === 5'b11111);
assign rom_instr_pt[197] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] , 
    rom_addr_l2[3] , rom_addr_l2[4] , 
    rom_addr_l2[6] }) === 5'b00001);
assign rom_instr_pt[198] =
    (({ rom_addr_l2[0] , rom_addr_l2[2] , 
    rom_addr_l2[3] , rom_addr_l2[4] , 
    rom_addr_l2[6] }) === 5'b00001);
assign rom_instr_pt[199] =
    (({ rom_addr_l2[1] , rom_addr_l2[3] , 
    rom_addr_l2[4] , rom_addr_l2[6]
     }) === 4'b0001);
assign rom_instr_pt[200] =
    (({ rom_addr_l2[0] , rom_addr_l2[3] , 
    rom_addr_l2[4] , rom_addr_l2[6]
     }) === 4'b0001);
assign rom_instr_pt[201] =
    (({ rom_addr_l2[0] , rom_addr_l2[2] , 
    rom_addr_l2[3] , rom_addr_l2[4] , 
    rom_addr_l2[6] }) === 5'b00011);
assign rom_instr_pt[202] =
    (({ rom_addr_l2[1] , rom_addr_l2[3] , 
    rom_addr_l2[4] , rom_addr_l2[6]
     }) === 4'b1111);
assign rom_instr_pt[203] =
    (({ rom_addr_l2[0] , rom_addr_l2[2] , 
    rom_addr_l2[4] , rom_addr_l2[6]
     }) === 4'b1111);
assign rom_instr_pt[204] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] , 
    rom_addr_l2[2] , rom_addr_l2[3] , 
    rom_addr_l2[6] }) === 5'b10001);
assign rom_instr_pt[205] =
    (({ rom_addr_l2[0] , rom_addr_l2[2] , 
    rom_addr_l2[3] , rom_addr_l2[6]
     }) === 4'b0001);
assign rom_instr_pt[206] =
    (({ rom_addr_l2[0] , rom_addr_l2[2] , 
    rom_addr_l2[3] , rom_addr_l2[6]
     }) === 4'b1111);
assign rom_instr_pt[207] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] , 
    rom_addr_l2[3] , rom_addr_l2[6]
     }) === 4'b0111);
assign rom_instr_pt[208] =
    (({ rom_addr_l2[2] , rom_addr_l2[6]
     }) === 2'b01);
assign rom_instr_pt[209] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] , 
    rom_addr_l2[2] , rom_addr_l2[3] , 
    rom_addr_l2[4] , rom_addr_l2[5]
     }) === 6'b011100);
assign rom_instr_pt[210] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] , 
    rom_addr_l2[4] , rom_addr_l2[5]
     }) === 4'b1010);
assign rom_instr_pt[211] =
    (({ rom_addr_l2[0] , rom_addr_l2[2] , 
    rom_addr_l2[3] , rom_addr_l2[5]
     }) === 4'b1000);
assign rom_instr_pt[212] =
    (({ rom_addr_l2[3] , rom_addr_l2[5]
     }) === 2'b00);
assign rom_instr_pt[213] =
    (({ rom_addr_l2[1] , rom_addr_l2[3] , 
    rom_addr_l2[5] }) === 3'b010);
assign rom_instr_pt[214] =
    (({ rom_addr_l2[1] , rom_addr_l2[3] , 
    rom_addr_l2[4] , rom_addr_l2[5]
     }) === 4'b1111);
assign rom_instr_pt[215] =
    (({ rom_addr_l2[0] , rom_addr_l2[2] , 
    rom_addr_l2[3] , rom_addr_l2[5]
     }) === 4'b0111);
assign rom_instr_pt[216] =
    (({ rom_addr_l2[0] , rom_addr_l2[2] , 
    rom_addr_l2[3] , rom_addr_l2[5]
     }) === 4'b1111);
assign rom_instr_pt[217] =
    (({ rom_addr_l2[0] , rom_addr_l2[2] , 
    rom_addr_l2[3] , rom_addr_l2[4]
     }) === 4'b1000);
assign rom_instr_pt[218] =
    (({ rom_addr_l2[3] , rom_addr_l2[4]
     }) === 2'b00);
assign rom_instr_pt[219] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] , 
    rom_addr_l2[3] , rom_addr_l2[4]
     }) === 4'b1001);
assign rom_instr_pt[220] =
    (({ rom_addr_l2[3] , rom_addr_l2[4]
     }) === 2'b11);
assign rom_instr_pt[221] =
    (({ rom_addr_l2[0] , rom_addr_l2[2] , 
    rom_addr_l2[4] }) === 3'b111);
assign rom_instr_pt[222] =
    (({ rom_addr_l2[1] , rom_addr_l2[4]
     }) === 2'b11);
assign rom_instr_pt[223] =
    (({ rom_addr_l2[0] , rom_addr_l2[2] , 
    rom_addr_l2[3] }) === 3'b111);
assign rom_instr_pt[224] =
    (({ rom_addr_l2[2] }) === 1'b0);
assign rom_instr_pt[225] =
    1'b1;
assign template[0] = 
    (rom_instr_pt[24] | rom_instr_pt[33]
     | rom_instr_pt[36] | rom_instr_pt[40]
     | rom_instr_pt[44] | rom_instr_pt[72]
     | rom_instr_pt[91] | rom_instr_pt[92]
     | rom_instr_pt[102] | rom_instr_pt[105]
     | rom_instr_pt[114] | rom_instr_pt[115]
     | rom_instr_pt[137] | rom_instr_pt[155]
     | rom_instr_pt[174] | rom_instr_pt[177]
     | rom_instr_pt[185] | rom_instr_pt[187]
     | rom_instr_pt[193] | rom_instr_pt[194]
     | rom_instr_pt[217]);
assign template[1] = 
    (rom_instr_pt[3] | rom_instr_pt[6]
     | rom_instr_pt[8] | rom_instr_pt[9]
     | rom_instr_pt[12] | rom_instr_pt[16]
     | rom_instr_pt[22] | rom_instr_pt[23]
     | rom_instr_pt[25] | rom_instr_pt[27]
     | rom_instr_pt[30] | rom_instr_pt[31]
     | rom_instr_pt[32] | rom_instr_pt[34]
     | rom_instr_pt[35] | rom_instr_pt[43]
     | rom_instr_pt[45] | rom_instr_pt[47]
     | rom_instr_pt[48] | rom_instr_pt[52]
     | rom_instr_pt[53] | rom_instr_pt[59]
     | rom_instr_pt[63] | rom_instr_pt[64]
     | rom_instr_pt[67] | rom_instr_pt[68]
     | rom_instr_pt[70] | rom_instr_pt[74]
     | rom_instr_pt[75] | rom_instr_pt[79]
     | rom_instr_pt[83] | rom_instr_pt[84]
     | rom_instr_pt[88] | rom_instr_pt[93]
     | rom_instr_pt[94] | rom_instr_pt[100]
     | rom_instr_pt[104] | rom_instr_pt[106]
     | rom_instr_pt[112] | rom_instr_pt[117]
     | rom_instr_pt[119] | rom_instr_pt[120]
     | rom_instr_pt[126] | rom_instr_pt[127]
     | rom_instr_pt[131] | rom_instr_pt[140]
     | rom_instr_pt[141] | rom_instr_pt[143]
     | rom_instr_pt[144] | rom_instr_pt[145]
     | rom_instr_pt[153] | rom_instr_pt[156]
     | rom_instr_pt[157] | rom_instr_pt[165]
     | rom_instr_pt[168] | rom_instr_pt[172]
     | rom_instr_pt[182] | rom_instr_pt[183]
     | rom_instr_pt[184] | rom_instr_pt[195]
     | rom_instr_pt[202] | rom_instr_pt[203]
     | rom_instr_pt[204] | rom_instr_pt[205]
     | rom_instr_pt[206] | rom_instr_pt[211]
     | rom_instr_pt[216]);
assign template[2] = 
    (rom_instr_pt[4] | rom_instr_pt[9]
     | rom_instr_pt[10] | rom_instr_pt[14]
     | rom_instr_pt[16] | rom_instr_pt[18]
     | rom_instr_pt[21] | rom_instr_pt[25]
     | rom_instr_pt[31] | rom_instr_pt[32]
     | rom_instr_pt[38] | rom_instr_pt[47]
     | rom_instr_pt[52] | rom_instr_pt[60]
     | rom_instr_pt[62] | rom_instr_pt[70]
     | rom_instr_pt[84] | rom_instr_pt[86]
     | rom_instr_pt[89] | rom_instr_pt[93]
     | rom_instr_pt[98] | rom_instr_pt[99]
     | rom_instr_pt[100] | rom_instr_pt[103]
     | rom_instr_pt[108] | rom_instr_pt[112]
     | rom_instr_pt[117] | rom_instr_pt[119]
     | rom_instr_pt[120] | rom_instr_pt[129]
     | rom_instr_pt[139] | rom_instr_pt[141]
     | rom_instr_pt[143] | rom_instr_pt[144]
     | rom_instr_pt[145] | rom_instr_pt[153]
     | rom_instr_pt[157] | rom_instr_pt[163]
     | rom_instr_pt[164] | rom_instr_pt[167]
     | rom_instr_pt[171] | rom_instr_pt[172]
     | rom_instr_pt[182] | rom_instr_pt[183]
     | rom_instr_pt[187] | rom_instr_pt[195]
     | rom_instr_pt[203] | rom_instr_pt[205]
     | rom_instr_pt[206] | rom_instr_pt[217]
    );
assign template[3] = 
    (rom_instr_pt[4] | rom_instr_pt[9]
     | rom_instr_pt[10] | rom_instr_pt[12]
     | rom_instr_pt[16] | rom_instr_pt[18]
     | rom_instr_pt[21] | rom_instr_pt[23]
     | rom_instr_pt[25] | rom_instr_pt[27]
     | rom_instr_pt[31] | rom_instr_pt[32]
     | rom_instr_pt[34] | rom_instr_pt[38]
     | rom_instr_pt[43] | rom_instr_pt[45]
     | rom_instr_pt[47] | rom_instr_pt[48]
     | rom_instr_pt[52] | rom_instr_pt[53]
     | rom_instr_pt[61] | rom_instr_pt[62]
     | rom_instr_pt[63] | rom_instr_pt[64]
     | rom_instr_pt[65] | rom_instr_pt[67]
     | rom_instr_pt[74] | rom_instr_pt[79]
     | rom_instr_pt[83] | rom_instr_pt[84]
     | rom_instr_pt[86] | rom_instr_pt[88]
     | rom_instr_pt[89] | rom_instr_pt[94]
     | rom_instr_pt[98] | rom_instr_pt[99]
     | rom_instr_pt[100] | rom_instr_pt[103]
     | rom_instr_pt[104] | rom_instr_pt[108]
     | rom_instr_pt[109] | rom_instr_pt[114]
     | rom_instr_pt[115] | rom_instr_pt[117]
     | rom_instr_pt[119] | rom_instr_pt[120]
     | rom_instr_pt[126] | rom_instr_pt[127]
     | rom_instr_pt[129] | rom_instr_pt[137]
     | rom_instr_pt[139] | rom_instr_pt[141]
     | rom_instr_pt[143] | rom_instr_pt[145]
     | rom_instr_pt[156] | rom_instr_pt[164]
     | rom_instr_pt[165] | rom_instr_pt[167]
     | rom_instr_pt[171] | rom_instr_pt[172]
     | rom_instr_pt[177] | rom_instr_pt[182]
     | rom_instr_pt[194] | rom_instr_pt[195]
     | rom_instr_pt[198] | rom_instr_pt[204]
     | rom_instr_pt[211] | rom_instr_pt[222]
    );
assign template[4] = 
    (rom_instr_pt[4] | rom_instr_pt[9]
     | rom_instr_pt[10] | rom_instr_pt[16]
     | rom_instr_pt[18] | rom_instr_pt[21]
     | rom_instr_pt[24] | rom_instr_pt[25]
     | rom_instr_pt[31] | rom_instr_pt[32]
     | rom_instr_pt[33] | rom_instr_pt[36]
     | rom_instr_pt[38] | rom_instr_pt[40]
     | rom_instr_pt[44] | rom_instr_pt[47]
     | rom_instr_pt[52] | rom_instr_pt[60]
     | rom_instr_pt[62] | rom_instr_pt[70]
     | rom_instr_pt[72] | rom_instr_pt[84]
     | rom_instr_pt[86] | rom_instr_pt[89]
     | rom_instr_pt[91] | rom_instr_pt[92]
     | rom_instr_pt[93] | rom_instr_pt[98]
     | rom_instr_pt[99] | rom_instr_pt[100]
     | rom_instr_pt[102] | rom_instr_pt[103]
     | rom_instr_pt[105] | rom_instr_pt[108]
     | rom_instr_pt[112] | rom_instr_pt[114]
     | rom_instr_pt[115] | rom_instr_pt[117]
     | rom_instr_pt[119] | rom_instr_pt[120]
     | rom_instr_pt[129] | rom_instr_pt[137]
     | rom_instr_pt[139] | rom_instr_pt[141]
     | rom_instr_pt[143] | rom_instr_pt[144]
     | rom_instr_pt[145] | rom_instr_pt[153]
     | rom_instr_pt[157] | rom_instr_pt[163]
     | rom_instr_pt[164] | rom_instr_pt[167]
     | rom_instr_pt[171] | rom_instr_pt[172]
     | rom_instr_pt[177] | rom_instr_pt[182]
     | rom_instr_pt[183] | rom_instr_pt[185]
     | rom_instr_pt[194] | rom_instr_pt[195]
     | rom_instr_pt[203] | rom_instr_pt[205]
     | rom_instr_pt[206] | rom_instr_pt[216]
     | rom_instr_pt[217]);
assign template[5] = 
    (rom_instr_pt[3] | rom_instr_pt[6]
     | rom_instr_pt[8] | rom_instr_pt[9]
     | rom_instr_pt[12] | rom_instr_pt[16]
     | rom_instr_pt[20] | rom_instr_pt[21]
     | rom_instr_pt[25] | rom_instr_pt[27]
     | rom_instr_pt[30] | rom_instr_pt[32]
     | rom_instr_pt[34] | rom_instr_pt[35]
     | rom_instr_pt[43] | rom_instr_pt[47]
     | rom_instr_pt[51] | rom_instr_pt[52]
     | rom_instr_pt[59] | rom_instr_pt[61]
     | rom_instr_pt[64] | rom_instr_pt[65]
     | rom_instr_pt[67] | rom_instr_pt[68]
     | rom_instr_pt[70] | rom_instr_pt[74]
     | rom_instr_pt[79] | rom_instr_pt[83]
     | rom_instr_pt[84] | rom_instr_pt[93]
     | rom_instr_pt[100] | rom_instr_pt[104]
     | rom_instr_pt[106] | rom_instr_pt[109]
     | rom_instr_pt[117] | rom_instr_pt[119]
     | rom_instr_pt[124] | rom_instr_pt[126]
     | rom_instr_pt[127] | rom_instr_pt[131]
     | rom_instr_pt[140] | rom_instr_pt[141]
     | rom_instr_pt[143] | rom_instr_pt[145]
     | rom_instr_pt[156] | rom_instr_pt[157]
     | rom_instr_pt[165] | rom_instr_pt[168]
     | rom_instr_pt[172] | rom_instr_pt[182]
     | rom_instr_pt[184] | rom_instr_pt[195]
     | rom_instr_pt[198] | rom_instr_pt[202]
     | rom_instr_pt[217]);
assign template[6] = 
    1'b0;
assign template[7] = 
    1'b0;
assign template[8] = 
    1'b0;
assign template[9] = 
    (rom_instr_pt[23] | rom_instr_pt[27]
     | rom_instr_pt[31] | rom_instr_pt[34]
     | rom_instr_pt[35] | rom_instr_pt[43]
     | rom_instr_pt[48] | rom_instr_pt[53]
     | rom_instr_pt[59] | rom_instr_pt[64]
     | rom_instr_pt[67] | rom_instr_pt[68]
     | rom_instr_pt[72] | rom_instr_pt[75]
     | rom_instr_pt[84] | rom_instr_pt[91]
     | rom_instr_pt[94] | rom_instr_pt[100]
     | rom_instr_pt[105] | rom_instr_pt[112]
     | rom_instr_pt[114] | rom_instr_pt[115]
     | rom_instr_pt[117] | rom_instr_pt[119]
     | rom_instr_pt[120] | rom_instr_pt[126]
     | rom_instr_pt[127] | rom_instr_pt[137]
     | rom_instr_pt[139] | rom_instr_pt[141]
     | rom_instr_pt[144] | rom_instr_pt[153]
     | rom_instr_pt[156] | rom_instr_pt[163]
     | rom_instr_pt[167] | rom_instr_pt[168]
     | rom_instr_pt[177] | rom_instr_pt[182]
     | rom_instr_pt[183] | rom_instr_pt[194]
     | rom_instr_pt[195]);
assign template[10] = 
    (rom_instr_pt[22] | rom_instr_pt[24]
     | rom_instr_pt[25] | rom_instr_pt[32]
     | rom_instr_pt[33] | rom_instr_pt[36]
     | rom_instr_pt[40] | rom_instr_pt[44]
     | rom_instr_pt[45] | rom_instr_pt[47]
     | rom_instr_pt[52] | rom_instr_pt[63]
     | rom_instr_pt[83] | rom_instr_pt[88]
     | rom_instr_pt[92] | rom_instr_pt[102]
     | rom_instr_pt[106] | rom_instr_pt[151]
     | rom_instr_pt[167] | rom_instr_pt[204]
     | rom_instr_pt[211]);
assign template[11] = 
    (rom_instr_pt[8] | rom_instr_pt[30]
     | rom_instr_pt[93] | rom_instr_pt[183]
    );
assign template[12] = 
    (rom_instr_pt[8] | rom_instr_pt[30]
    );
assign template[13] = 
    1'b0;
assign template[14] = 
    (rom_instr_pt[12] | rom_instr_pt[27]
     | rom_instr_pt[31] | rom_instr_pt[34]
     | rom_instr_pt[43] | rom_instr_pt[45]
     | rom_instr_pt[53] | rom_instr_pt[59]
     | rom_instr_pt[63] | rom_instr_pt[64]
     | rom_instr_pt[67] | rom_instr_pt[70]
     | rom_instr_pt[75] | rom_instr_pt[79]
     | rom_instr_pt[83] | rom_instr_pt[88]
     | rom_instr_pt[93] | rom_instr_pt[94]
     | rom_instr_pt[104] | rom_instr_pt[117]
     | rom_instr_pt[120] | rom_instr_pt[126]
     | rom_instr_pt[127] | rom_instr_pt[131]
     | rom_instr_pt[156] | rom_instr_pt[165]
     | rom_instr_pt[168] | rom_instr_pt[204]
     | rom_instr_pt[211]);
assign template[15] = 
    (rom_instr_pt[3] | rom_instr_pt[23]
     | rom_instr_pt[48] | rom_instr_pt[172]
     | rom_instr_pt[175] | rom_instr_pt[202]
    );
assign template[16] = 
    (rom_instr_pt[4] | rom_instr_pt[34]
     | rom_instr_pt[51] | rom_instr_pt[53]
     | rom_instr_pt[63] | rom_instr_pt[75]
     | rom_instr_pt[94] | rom_instr_pt[120]
     | rom_instr_pt[151] | rom_instr_pt[165]
     | rom_instr_pt[204]);
assign template[17] = 
    (rom_instr_pt[4] | rom_instr_pt[12]
     | rom_instr_pt[27] | rom_instr_pt[31]
     | rom_instr_pt[34] | rom_instr_pt[43]
     | rom_instr_pt[45] | rom_instr_pt[59]
     | rom_instr_pt[63] | rom_instr_pt[64]
     | rom_instr_pt[67] | rom_instr_pt[75]
     | rom_instr_pt[79] | rom_instr_pt[83]
     | rom_instr_pt[88] | rom_instr_pt[104]
     | rom_instr_pt[120] | rom_instr_pt[126]
     | rom_instr_pt[127] | rom_instr_pt[131]
     | rom_instr_pt[151] | rom_instr_pt[156]
     | rom_instr_pt[168] | rom_instr_pt[204]
    );
assign template[18] = 
    (rom_instr_pt[4] | rom_instr_pt[124]
     | rom_instr_pt[151]);
assign template[19] = 
    (rom_instr_pt[4] | rom_instr_pt[145]
     | rom_instr_pt[151]);
assign template[20] = 
    (rom_instr_pt[4] | rom_instr_pt[56]
     | rom_instr_pt[70] | rom_instr_pt[84]
     | rom_instr_pt[117] | rom_instr_pt[137]
     | rom_instr_pt[151] | rom_instr_pt[175]
    );
assign template[21] = 
    (rom_instr_pt[4] | rom_instr_pt[22]
     | rom_instr_pt[23] | rom_instr_pt[43]
     | rom_instr_pt[45] | rom_instr_pt[48]
     | rom_instr_pt[53] | rom_instr_pt[88]
     | rom_instr_pt[94] | rom_instr_pt[109]
     | rom_instr_pt[145] | rom_instr_pt[151]
    );
assign template[22] = 
    (rom_instr_pt[3] | rom_instr_pt[4]
     | rom_instr_pt[23] | rom_instr_pt[48]
     | rom_instr_pt[61] | rom_instr_pt[65]
     | rom_instr_pt[70] | rom_instr_pt[84]
     | rom_instr_pt[109] | rom_instr_pt[117]
     | rom_instr_pt[140] | rom_instr_pt[143]
     | rom_instr_pt[151] | rom_instr_pt[157]
     | rom_instr_pt[172] | rom_instr_pt[184]
     | rom_instr_pt[198] | rom_instr_pt[202]
    );
assign template[23] = 
    (rom_instr_pt[4] | rom_instr_pt[22]
     | rom_instr_pt[30] | rom_instr_pt[35]
     | rom_instr_pt[51] | rom_instr_pt[68]
     | rom_instr_pt[84] | rom_instr_pt[93]
     | rom_instr_pt[100] | rom_instr_pt[109]
     | rom_instr_pt[117] | rom_instr_pt[119]
     | rom_instr_pt[124] | rom_instr_pt[141]
     | rom_instr_pt[151] | rom_instr_pt[157]
     | rom_instr_pt[182] | rom_instr_pt[184]
     | rom_instr_pt[195] | rom_instr_pt[202]
    );
assign template[24] = 
    (rom_instr_pt[3] | rom_instr_pt[4]
     | rom_instr_pt[22] | rom_instr_pt[25]
     | rom_instr_pt[32] | rom_instr_pt[35]
     | rom_instr_pt[47] | rom_instr_pt[52]
     | rom_instr_pt[68] | rom_instr_pt[74]
     | rom_instr_pt[100] | rom_instr_pt[106]
     | rom_instr_pt[119] | rom_instr_pt[139]
     | rom_instr_pt[141] | rom_instr_pt[145]
     | rom_instr_pt[151] | rom_instr_pt[182]
     | rom_instr_pt[195]);
assign template[25] = 
    (rom_instr_pt[4] | rom_instr_pt[20]
     | rom_instr_pt[21] | rom_instr_pt[60]
     | rom_instr_pt[70] | rom_instr_pt[84]
     | rom_instr_pt[117] | rom_instr_pt[145]
     | rom_instr_pt[151] | rom_instr_pt[157]
     | rom_instr_pt[184]);
assign template[26] = 
    (rom_instr_pt[3] | rom_instr_pt[4]
     | rom_instr_pt[6] | rom_instr_pt[8]
     | rom_instr_pt[9] | rom_instr_pt[12]
     | rom_instr_pt[16] | rom_instr_pt[22]
     | rom_instr_pt[23] | rom_instr_pt[25]
     | rom_instr_pt[27] | rom_instr_pt[30]
     | rom_instr_pt[32] | rom_instr_pt[34]
     | rom_instr_pt[35] | rom_instr_pt[43]
     | rom_instr_pt[45] | rom_instr_pt[47]
     | rom_instr_pt[48] | rom_instr_pt[51]
     | rom_instr_pt[52] | rom_instr_pt[53]
     | rom_instr_pt[59] | rom_instr_pt[64]
     | rom_instr_pt[67] | rom_instr_pt[68]
     | rom_instr_pt[70] | rom_instr_pt[74]
     | rom_instr_pt[79] | rom_instr_pt[83]
     | rom_instr_pt[84] | rom_instr_pt[88]
     | rom_instr_pt[93] | rom_instr_pt[94]
     | rom_instr_pt[100] | rom_instr_pt[104]
     | rom_instr_pt[106] | rom_instr_pt[109]
     | rom_instr_pt[117] | rom_instr_pt[119]
     | rom_instr_pt[124] | rom_instr_pt[126]
     | rom_instr_pt[127] | rom_instr_pt[131]
     | rom_instr_pt[141] | rom_instr_pt[145]
     | rom_instr_pt[151] | rom_instr_pt[156]
     | rom_instr_pt[157] | rom_instr_pt[168]
     | rom_instr_pt[182] | rom_instr_pt[184]
     | rom_instr_pt[195] | rom_instr_pt[202]
     | rom_instr_pt[211]);
assign template[27] = 
    (rom_instr_pt[4] | rom_instr_pt[6]
     | rom_instr_pt[9] | rom_instr_pt[12]
     | rom_instr_pt[16] | rom_instr_pt[20]
     | rom_instr_pt[21] | rom_instr_pt[23]
     | rom_instr_pt[27] | rom_instr_pt[34]
     | rom_instr_pt[48] | rom_instr_pt[59]
     | rom_instr_pt[60] | rom_instr_pt[61]
     | rom_instr_pt[64] | rom_instr_pt[65]
     | rom_instr_pt[79] | rom_instr_pt[83]
     | rom_instr_pt[84] | rom_instr_pt[104]
     | rom_instr_pt[109] | rom_instr_pt[117]
     | rom_instr_pt[126] | rom_instr_pt[127]
     | rom_instr_pt[130] | rom_instr_pt[131]
     | rom_instr_pt[140] | rom_instr_pt[143]
     | rom_instr_pt[145] | rom_instr_pt[151]
     | rom_instr_pt[157] | rom_instr_pt[168]
     | rom_instr_pt[172] | rom_instr_pt[184]
     | rom_instr_pt[198] | rom_instr_pt[209]
    );
assign template[28] = 
    (rom_instr_pt[4] | rom_instr_pt[6]
     | rom_instr_pt[9] | rom_instr_pt[12]
     | rom_instr_pt[16] | rom_instr_pt[20]
     | rom_instr_pt[21] | rom_instr_pt[23]
     | rom_instr_pt[25] | rom_instr_pt[27]
     | rom_instr_pt[32] | rom_instr_pt[34]
     | rom_instr_pt[35] | rom_instr_pt[43]
     | rom_instr_pt[45] | rom_instr_pt[47]
     | rom_instr_pt[48] | rom_instr_pt[52]
     | rom_instr_pt[53] | rom_instr_pt[59]
     | rom_instr_pt[60] | rom_instr_pt[63]
     | rom_instr_pt[64] | rom_instr_pt[67]
     | rom_instr_pt[68] | rom_instr_pt[70]
     | rom_instr_pt[74] | rom_instr_pt[79]
     | rom_instr_pt[83] | rom_instr_pt[84]
     | rom_instr_pt[88] | rom_instr_pt[94]
     | rom_instr_pt[100] | rom_instr_pt[104]
     | rom_instr_pt[106] | rom_instr_pt[117]
     | rom_instr_pt[119] | rom_instr_pt[126]
     | rom_instr_pt[127] | rom_instr_pt[131]
     | rom_instr_pt[141] | rom_instr_pt[145]
     | rom_instr_pt[151] | rom_instr_pt[156]
     | rom_instr_pt[157] | rom_instr_pt[165]
     | rom_instr_pt[168] | rom_instr_pt[182]
     | rom_instr_pt[184] | rom_instr_pt[195]
     | rom_instr_pt[204]);
assign template[29] = 
    (rom_instr_pt[3] | rom_instr_pt[4]
     | rom_instr_pt[8] | rom_instr_pt[12]
     | rom_instr_pt[20] | rom_instr_pt[21]
     | rom_instr_pt[23] | rom_instr_pt[25]
     | rom_instr_pt[27] | rom_instr_pt[32]
     | rom_instr_pt[34] | rom_instr_pt[35]
     | rom_instr_pt[43] | rom_instr_pt[45]
     | rom_instr_pt[47] | rom_instr_pt[48]
     | rom_instr_pt[52] | rom_instr_pt[53]
     | rom_instr_pt[59] | rom_instr_pt[61]
     | rom_instr_pt[63] | rom_instr_pt[64]
     | rom_instr_pt[65] | rom_instr_pt[67]
     | rom_instr_pt[68] | rom_instr_pt[74]
     | rom_instr_pt[79] | rom_instr_pt[83]
     | rom_instr_pt[86] | rom_instr_pt[88]
     | rom_instr_pt[94] | rom_instr_pt[100]
     | rom_instr_pt[104] | rom_instr_pt[106]
     | rom_instr_pt[109] | rom_instr_pt[119]
     | rom_instr_pt[126] | rom_instr_pt[127]
     | rom_instr_pt[131] | rom_instr_pt[139]
     | rom_instr_pt[141] | rom_instr_pt[143]
     | rom_instr_pt[145] | rom_instr_pt[151]
     | rom_instr_pt[156] | rom_instr_pt[165]
     | rom_instr_pt[168] | rom_instr_pt[172]
     | rom_instr_pt[182] | rom_instr_pt[195]
     | rom_instr_pt[198] | rom_instr_pt[204]
    );
assign template[30] = 
    (rom_instr_pt[4] | rom_instr_pt[12]
     | rom_instr_pt[15] | rom_instr_pt[20]
     | rom_instr_pt[23] | rom_instr_pt[24]
     | rom_instr_pt[25] | rom_instr_pt[27]
     | rom_instr_pt[32] | rom_instr_pt[34]
     | rom_instr_pt[35] | rom_instr_pt[43]
     | rom_instr_pt[45] | rom_instr_pt[47]
     | rom_instr_pt[48] | rom_instr_pt[52]
     | rom_instr_pt[53] | rom_instr_pt[59]
     | rom_instr_pt[63] | rom_instr_pt[64]
     | rom_instr_pt[67] | rom_instr_pt[68]
     | rom_instr_pt[74] | rom_instr_pt[75]
     | rom_instr_pt[79] | rom_instr_pt[83]
     | rom_instr_pt[88] | rom_instr_pt[94]
     | rom_instr_pt[100] | rom_instr_pt[102]
     | rom_instr_pt[104] | rom_instr_pt[106]
     | rom_instr_pt[119] | rom_instr_pt[120]
     | rom_instr_pt[126] | rom_instr_pt[127]
     | rom_instr_pt[131] | rom_instr_pt[139]
     | rom_instr_pt[141] | rom_instr_pt[145]
     | rom_instr_pt[156] | rom_instr_pt[165]
     | rom_instr_pt[168] | rom_instr_pt[182]
     | rom_instr_pt[195] | rom_instr_pt[204]
    );
assign template[31] = 
    (rom_instr_pt[14] | rom_instr_pt[24]
     | rom_instr_pt[33] | rom_instr_pt[38]
     | rom_instr_pt[62] | rom_instr_pt[77]
     | rom_instr_pt[89] | rom_instr_pt[91]
     | rom_instr_pt[98] | rom_instr_pt[99]
     | rom_instr_pt[103] | rom_instr_pt[108]
     | rom_instr_pt[122] | rom_instr_pt[170]
    );
assign ucode_end = 
    (rom_instr_pt[107] | rom_instr_pt[139]
     | rom_instr_pt[146] | rom_instr_pt[152]
     | rom_instr_pt[154] | rom_instr_pt[159]
     | rom_instr_pt[160] | rom_instr_pt[172]
     | rom_instr_pt[176] | rom_instr_pt[205]
     | rom_instr_pt[209]);
assign ucode_end_early = 
    (rom_instr_pt[87] | rom_instr_pt[111]
     | rom_instr_pt[125] | rom_instr_pt[207]
    );
assign loop_begin = 
    (rom_instr_pt[36] | rom_instr_pt[62]
     | rom_instr_pt[66] | rom_instr_pt[68]
     | rom_instr_pt[71] | rom_instr_pt[80]
     | rom_instr_pt[81] | rom_instr_pt[96]
     | rom_instr_pt[105] | rom_instr_pt[106]
     | rom_instr_pt[121] | rom_instr_pt[123]
     | rom_instr_pt[132] | rom_instr_pt[133]
     | rom_instr_pt[135]);
assign loop_end = 
    (rom_instr_pt[55] | rom_instr_pt[87]
     | rom_instr_pt[158] | rom_instr_pt[199]
     | rom_instr_pt[200] | rom_instr_pt[208]
     | rom_instr_pt[209]);
assign count_src[0] = 
    (rom_instr_pt[189] | rom_instr_pt[212]
     | rom_instr_pt[218] | rom_instr_pt[224]
    );
assign count_src[1] = 
    (rom_instr_pt[161] | rom_instr_pt[218]
     | rom_instr_pt[220] | rom_instr_pt[224]
    );
assign count_src[2] = 
    (rom_instr_pt[188] | rom_instr_pt[213]
     | rom_instr_pt[218] | rom_instr_pt[224]
    );
assign ext_rt = 
    (rom_instr_pt[1] | rom_instr_pt[4]
     | rom_instr_pt[6] | rom_instr_pt[9]
     | rom_instr_pt[11] | rom_instr_pt[12]
     | rom_instr_pt[13] | rom_instr_pt[19]
     | rom_instr_pt[21] | rom_instr_pt[23]
     | rom_instr_pt[28] | rom_instr_pt[32]
     | rom_instr_pt[37] | rom_instr_pt[41]
     | rom_instr_pt[42] | rom_instr_pt[43]
     | rom_instr_pt[47] | rom_instr_pt[48]
     | rom_instr_pt[49] | rom_instr_pt[52]
     | rom_instr_pt[54] | rom_instr_pt[58]
     | rom_instr_pt[61] | rom_instr_pt[63]
     | rom_instr_pt[65] | rom_instr_pt[67]
     | rom_instr_pt[69] | rom_instr_pt[76]
     | rom_instr_pt[82] | rom_instr_pt[97]
     | rom_instr_pt[113] | rom_instr_pt[118]
     | rom_instr_pt[120] | rom_instr_pt[128]
     | rom_instr_pt[134] | rom_instr_pt[142]
     | rom_instr_pt[147] | rom_instr_pt[166]
     | rom_instr_pt[173] | rom_instr_pt[181]
     | rom_instr_pt[186] | rom_instr_pt[204]
     | rom_instr_pt[210] | rom_instr_pt[215]
     | rom_instr_pt[219]);
assign ext_s1 = 
    (rom_instr_pt[23] | rom_instr_pt[28]
     | rom_instr_pt[41] | rom_instr_pt[42]
     | rom_instr_pt[48] | rom_instr_pt[50]
     | rom_instr_pt[54] | rom_instr_pt[57]
     | rom_instr_pt[58] | rom_instr_pt[63]
     | rom_instr_pt[67] | rom_instr_pt[69]
     | rom_instr_pt[76] | rom_instr_pt[82]
     | rom_instr_pt[90] | rom_instr_pt[101]
     | rom_instr_pt[113] | rom_instr_pt[115]
     | rom_instr_pt[116] | rom_instr_pt[118]
     | rom_instr_pt[134] | rom_instr_pt[147]
     | rom_instr_pt[148] | rom_instr_pt[149]
     | rom_instr_pt[155] | rom_instr_pt[162]
     | rom_instr_pt[166] | rom_instr_pt[169]
     | rom_instr_pt[172] | rom_instr_pt[173]
     | rom_instr_pt[178] | rom_instr_pt[179]
     | rom_instr_pt[181] | rom_instr_pt[201]
     | rom_instr_pt[204] | rom_instr_pt[210]
     | rom_instr_pt[219]);
assign ext_s2 = 
    (rom_instr_pt[23] | rom_instr_pt[32]
     | rom_instr_pt[47] | rom_instr_pt[48]
     | rom_instr_pt[52] | rom_instr_pt[54]
     | rom_instr_pt[63] | rom_instr_pt[85]
     | rom_instr_pt[90] | rom_instr_pt[95]
     | rom_instr_pt[145] | rom_instr_pt[148]
     | rom_instr_pt[172] | rom_instr_pt[181]
     | rom_instr_pt[197] | rom_instr_pt[204]
     | rom_instr_pt[210] | rom_instr_pt[214]
    );
assign ext_s3 = 
    (rom_instr_pt[46] | rom_instr_pt[58]
     | rom_instr_pt[68] | rom_instr_pt[115]
     | rom_instr_pt[116] | rom_instr_pt[119]
     | rom_instr_pt[134] | rom_instr_pt[147]
     | rom_instr_pt[149] | rom_instr_pt[178]
     | rom_instr_pt[215]);
assign sel0_5 = 
    (rom_instr_pt[148]);
assign sel6_10[0] = 
    (rom_instr_pt[6] | rom_instr_pt[9]
     | rom_instr_pt[19] | rom_instr_pt[136]
     | rom_instr_pt[146] | rom_instr_pt[150]
     | rom_instr_pt[172] | rom_instr_pt[198]
    );
assign sel6_10[1] = 
    (rom_instr_pt[6] | rom_instr_pt[9]
     | rom_instr_pt[11] | rom_instr_pt[12]
     | rom_instr_pt[19] | rom_instr_pt[37]
     | rom_instr_pt[73] | rom_instr_pt[79]
     | rom_instr_pt[97] | rom_instr_pt[104]
     | rom_instr_pt[145] | rom_instr_pt[148]
     | rom_instr_pt[155] | rom_instr_pt[174]
     | rom_instr_pt[191] | rom_instr_pt[193]
     | rom_instr_pt[214]);
assign sel11_15[0] = 
    (rom_instr_pt[85] | rom_instr_pt[110]
     | rom_instr_pt[153] | rom_instr_pt[157]
     | rom_instr_pt[179] | rom_instr_pt[180]
     | rom_instr_pt[196]);
assign sel11_15[1] = 
    (rom_instr_pt[1] | rom_instr_pt[4]
     | rom_instr_pt[7] | rom_instr_pt[13]
     | rom_instr_pt[32] | rom_instr_pt[46]
     | rom_instr_pt[47] | rom_instr_pt[49]
     | rom_instr_pt[52] | rom_instr_pt[85]
     | rom_instr_pt[110] | rom_instr_pt[128]
     | rom_instr_pt[136] | rom_instr_pt[142]
     | rom_instr_pt[146] | rom_instr_pt[150]
     | rom_instr_pt[153] | rom_instr_pt[157]
     | rom_instr_pt[179] | rom_instr_pt[180]
     | rom_instr_pt[196] | rom_instr_pt[197]
     | rom_instr_pt[201] | rom_instr_pt[221]
     | rom_instr_pt[223]);
assign sel16_20[0] = 
    (rom_instr_pt[17] | rom_instr_pt[20]
     | rom_instr_pt[21]);
assign sel16_20[1] = 
    (rom_instr_pt[1] | rom_instr_pt[2]
     | rom_instr_pt[6] | rom_instr_pt[9]
     | rom_instr_pt[19] | rom_instr_pt[26]
     | rom_instr_pt[29] | rom_instr_pt[35]
     | rom_instr_pt[39] | rom_instr_pt[42]
     | rom_instr_pt[46] | rom_instr_pt[57]
     | rom_instr_pt[61] | rom_instr_pt[65]
     | rom_instr_pt[68] | rom_instr_pt[74]
     | rom_instr_pt[101] | rom_instr_pt[106]
     | rom_instr_pt[115] | rom_instr_pt[116]
     | rom_instr_pt[119] | rom_instr_pt[136]
     | rom_instr_pt[146] | rom_instr_pt[149]
     | rom_instr_pt[150] | rom_instr_pt[190]
     | rom_instr_pt[191] | rom_instr_pt[193]
     | rom_instr_pt[195]);
assign sel21_25[0] = 
    1'b0;
assign sel21_25[1] = 
    (rom_instr_pt[1] | rom_instr_pt[2]
     | rom_instr_pt[29] | rom_instr_pt[39]
     | rom_instr_pt[42] | rom_instr_pt[115]
     | rom_instr_pt[136] | rom_instr_pt[138]
     | rom_instr_pt[191] | rom_instr_pt[193]
    );
assign sel26_30 = 
    (rom_instr_pt[1] | rom_instr_pt[2]
     | rom_instr_pt[29] | rom_instr_pt[39]
     | rom_instr_pt[42] | rom_instr_pt[115]
     | rom_instr_pt[136] | rom_instr_pt[138]
     | rom_instr_pt[191] | rom_instr_pt[193]
    );
assign sel31 = 
    (rom_instr_pt[2] | rom_instr_pt[5]
     | rom_instr_pt[29] | rom_instr_pt[39]
     | rom_instr_pt[42] | rom_instr_pt[136]
     | rom_instr_pt[148] | rom_instr_pt[149]
     | rom_instr_pt[191] | rom_instr_pt[192]
    );
assign cr_bf2fxm = 
    1'b0;
assign skip_cond = 
    (rom_instr_pt[23] | rom_instr_pt[43]
     | rom_instr_pt[48] | rom_instr_pt[54]
     | rom_instr_pt[63] | rom_instr_pt[78]
     | rom_instr_pt[95] | rom_instr_pt[113]
     | rom_instr_pt[118] | rom_instr_pt[120]
     | rom_instr_pt[204]);
assign skip_zero = 
    (rom_instr_pt[67] | rom_instr_pt[155]
     | rom_instr_pt[166] | rom_instr_pt[186]
     | rom_instr_pt[215]);
assign skip_nop = 
    1'b0;
assign loop_addr[0] = 
    1'b0;
assign loop_addr[1] = 
    1'b0;
assign loop_addr[2] = 
    1'b0;
assign loop_addr[3] = 
    1'b0;
assign loop_addr[4] = 
    1'b0;
assign loop_addr[5] = 
    1'b0;
assign loop_addr[6] = 
    1'b0;
assign loop_addr[7] = 
    1'b0;
assign loop_addr[8] = 
    1'b0;
assign loop_addr[9] = 
    1'b0;
assign loop_init[0] = 
    (rom_instr_pt[69] | rom_instr_pt[76]
     | rom_instr_pt[115] | rom_instr_pt[116]
     | rom_instr_pt[120]);
assign loop_init[1] = 
    (rom_instr_pt[225]);
assign loop_init[2] = 
    (rom_instr_pt[78]);
assign ep = 
    (rom_instr_pt[32] | rom_instr_pt[46]
     | rom_instr_pt[47] | rom_instr_pt[116]
     | rom_instr_pt[149] | rom_instr_pt[195]
    );





   assign rom_addr_d = rom_addr;

   assign rom_data = {template, ucode_end, ucode_end_early, loop_begin, loop_end, count_src, ext_rt, ext_s1, ext_s2, ext_s3, sel0_5, sel6_10, sel11_15, sel16_20, sel21_25, sel26_30, sel31, cr_bf2fxm, skip_cond, skip_zero, skip_nop, loop_addr, loop_init, ep};


   tri_rlmreg_p #(.WIDTH(10), .INIT(0), .NEEDS_SRESET(0)) rom_addr_latch(
      .vd(vdd),
      .gd(gnd),
      .nclk(nclk),
      .act(rom_act),
      .thold_b(pc_iu_func_sl_thold_0_b),
      .sg(pc_iu_sg_0),
      .force_t(force_t),
      .delay_lclkr(delay_lclkr),
      .mpw1_b(mpw1_b),
      .mpw2_b(mpw2_b),
      .d_mode(d_mode),
      .scin(siv[rom_addr_offset:rom_addr_offset + 10 - 1]),
      .scout(sov[rom_addr_offset:rom_addr_offset + 10 - 1]),
      .din(rom_addr_d),
      .dout(rom_addr_l2)
   );

   assign siv[0:scan_right] = {sov[1:scan_right], scan_in};
   assign scan_out = sov[0];

endmodule

