// © IBM Corp. 2020
// This softcore is licensed under and subject to the terms of the CC-BY 4.0
// license (https://creativecommons.org/licenses/by/4.0/legalcode). 
// Additional rights, including the right to physically implement a softcore 
// that is compliant with the required sections of the Power ISA 
// Specification, will be available at no cost via the OpenPOWER Foundation. 
// This README will be updated with additional information when OpenPOWER's 
// license is available.

`timescale 1 ns / 1 ns





module fu_gst_loa(
   a,
   shamt
);
   `include "tri_a2o.vh"
   
   
   input [1:19] a;
   
   output [0:4] shamt;
   
   
   wire         unused;
   
   assign unused = a[19];
   
   
   
   
   
   assign shamt[0] = ((~a[01]) & (~a[02]) & (~a[03]) & (~a[04]) & (~a[05]) & (~a[06]) & (~a[07]) & (~a[08]) & (~a[09]) & (~a[10]) & (~a[11]) & (~a[12]) & (~a[13]) & (~a[14]) & (~a[15]) & a[19]) | ((~a[01]) & (~a[02]) & (~a[03]) & (~a[04]) & (~a[05]) & (~a[06]) & (~a[07]) & (~a[08]) & (~a[09]) & (~a[10]) & (~a[11]) & (~a[12]) & (~a[13]) & (~a[14]) & (~a[15]) & a[18]) | ((~a[01]) & (~a[02]) & (~a[03]) & (~a[04]) & (~a[05]) & (~a[06]) & (~a[07]) & (~a[08]) & (~a[09]) & (~a[10]) & (~a[11]) & (~a[12]) & (~a[13]) & (~a[14]) & (~a[15]) & a[17]) | ((~a[01]) & (~a[02]) & (~a[03]) & (~a[04]) & (~a[05]) & (~a[06]) & (~a[07]) & (~a[08]) & (~a[09]) & (~a[10]) & (~a[11]) & (~a[12]) & (~a[13]) & (~a[14]) & (~a[15]) & a[16]);
   
   assign shamt[1] = ((~a[01]) & (~a[02]) & (~a[03]) & (~a[04]) & (~a[05]) & (~a[06]) & (~a[07]) & a[15]) | ((~a[01]) & (~a[02]) & (~a[03]) & (~a[04]) & (~a[05]) & (~a[06]) & (~a[07]) & a[14]) | ((~a[01]) & (~a[02]) & (~a[03]) & (~a[04]) & (~a[05]) & (~a[06]) & (~a[07]) & a[13]) | ((~a[01]) & (~a[02]) & (~a[03]) & (~a[04]) & (~a[05]) & (~a[06]) & (~a[07]) & a[12]) | ((~a[01]) & (~a[02]) & (~a[03]) & (~a[04]) & (~a[05]) & (~a[06]) & (~a[07]) & a[11]) | ((~a[01]) & (~a[02]) & (~a[03]) & (~a[04]) & (~a[05]) & (~a[06]) & (~a[07]) & a[10]) | ((~a[01]) & (~a[02]) & (~a[03]) & (~a[04]) & (~a[05]) & (~a[06]) & (~a[07]) & a[09]) | ((~a[01]) & (~a[02]) & (~a[03]) & (~a[04]) & (~a[05]) & (~a[06]) & (~a[07]) & a[08]);
   
   assign shamt[2] = ((~a[01]) & (~a[02]) & (~a[03]) & (~a[08]) & (~a[09]) & (~a[10]) & (~a[11]) & a[15]) | ((~a[01]) & (~a[02]) & (~a[03]) & (~a[08]) & (~a[09]) & (~a[10]) & (~a[11]) & a[14]) | ((~a[01]) & (~a[02]) & (~a[03]) & (~a[08]) & (~a[09]) & (~a[10]) & (~a[11]) & a[13]) | ((~a[01]) & (~a[02]) & (~a[03]) & (~a[08]) & (~a[09]) & (~a[10]) & (~a[11]) & a[12]) | ((~a[01]) & (~a[02]) & (~a[03]) & a[07]) | ((~a[01]) & (~a[02]) & (~a[03]) & a[06]) | ((~a[01]) & (~a[02]) & (~a[03]) & a[05]) | ((~a[01]) & (~a[02]) & (~a[03]) & a[04]);
   
   assign shamt[3] = ((~a[01]) & (~a[04]) & (~a[05]) & (~a[08]) & (~a[09]) & (~a[12]) & (~a[13]) & (~a[16]) & (~a[17]) & a[19]) | ((~a[01]) & (~a[04]) & (~a[05]) & (~a[08]) & (~a[09]) & (~a[12]) & (~a[13]) & (~a[16]) & (~a[17]) & a[18]) | ((~a[01]) & (~a[04]) & (~a[05]) & (~a[08]) & (~a[09]) & (~a[12]) & (~a[13]) & a[15]) | ((~a[01]) & (~a[04]) & (~a[05]) & (~a[08]) & (~a[09]) & (~a[12]) & (~a[13]) & a[14]) | ((~a[01]) & (~a[04]) & (~a[05]) & (~a[08]) & (~a[09]) & a[11]) | ((~a[01]) & (~a[04]) & (~a[05]) & (~a[08]) & (~a[09]) & a[10]) | ((~a[01]) & (~a[04]) & (~a[05]) & a[07]) | ((~a[01]) & (~a[04]) & (~a[05]) & a[06]) | ((~a[01]) & a[03]) | ((~a[01]) & a[02]);
   
   assign shamt[4] = ((~a[02]) & (~a[04]) & (~a[06]) & (~a[08]) & (~a[10]) & (~a[12]) & (~a[14]) & (~a[16]) & (~a[18]) & a[19]) | ((~a[02]) & (~a[04]) & (~a[06]) & (~a[08]) & (~a[10]) & (~a[12]) & (~a[14]) & (~a[16]) & a[17]) | ((~a[02]) & (~a[04]) & (~a[06]) & (~a[08]) & (~a[10]) & (~a[12]) & (~a[14]) & a[15]) | ((~a[02]) & (~a[04]) & (~a[06]) & (~a[08]) & (~a[10]) & (~a[12]) & a[13]) | ((~a[02]) & (~a[04]) & (~a[06]) & (~a[08]) & (~a[10]) & a[11]) | ((~a[02]) & (~a[04]) & (~a[06]) & (~a[08]) & a[09]) | ((~a[02]) & (~a[04]) & (~a[06]) & a[07]) | ((~a[02]) & (~a[04]) & a[05]) | ((~a[02]) & a[03]) | (a[01]);
   
endmodule
