// © IBM Corp. 2020
// This softcore is licensed under and subject to the terms of the CC-BY 4.0
// license (https://creativecommons.org/licenses/by/4.0/legalcode). 
// Additional rights, including the right to physically implement a softcore 
// that is compliant with the required sections of the Power ISA 
// Specification, will be available at no cost via the OpenPOWER Foundation. 
// This README will be updated with additional information when OpenPOWER's 
// license is available.

//********************************************************************
//*
//* TITLE: IU Microcode Code
//*
//* NAME: iuq_uc_rom_odd.v
//*
//*********************************************************************

`include "tri_a2o.vh"


module iuq_uc_rom_odd(
   vdd,
   gnd,
   nclk,
   pc_iu_func_sl_thold_0_b,
   pc_iu_sg_0,
   force_t,
   d_mode,
   delay_lclkr,
   mpw1_b,
   mpw2_b,
   scan_in,
   scan_out,
   rom_act,
   rom_addr,
   rom_data
);
   //parameter                ucode_width = 72;


   inout                    vdd;

   inout                    gnd;

    (* pin_data ="PIN_FUNCTION=/G_CLK/" *)
   input [0:`NCLK_WIDTH-1]  nclk;
   input                    pc_iu_func_sl_thold_0_b;
   input                    pc_iu_sg_0;
   input                    force_t;
   input                    d_mode;
   input                    delay_lclkr;
   input                    mpw1_b;
   input                    mpw2_b;
   input                    scan_in;
   output                   scan_out;

   input                    rom_act;
   input [0:9]              rom_addr;
   output [0:71]            rom_data;

   //@@  Signal Declarations
   wire [1:200]             rom_instr_pt;
   wire [0:2]               count_src;
   wire                     cr_bf2fxm;
   wire                     ep;
   wire                     ext_rt;
   wire                     ext_s1;
   wire                     ext_s2;
   wire                     ext_s3;
   wire [0:9]               loop_addr;
   wire                     loop_begin;
   wire                     loop_end;
   wire [0:2]               loop_init;
   wire                     sel0_5;
   wire [0:1]               sel11_15;
   wire [0:1]               sel16_20;
   wire [0:1]               sel21_25;
   wire                     sel26_30;
   wire                     sel31;
   wire [0:1]               sel6_10;
   wire                     skip_cond;
   wire                     skip_nop;
   wire                     skip_zero;
   wire [0:31]              template;
   wire                     ucode_end;
   wire                     ucode_end_early;

   parameter                rom_addr_offset = 0;
   parameter                scan_right = rom_addr_offset + 10 - 1;

   // Latches
   wire [0:9]               rom_addr_d;
   wire [0:9]               rom_addr_l2;
   wire [0:scan_right]      siv;
   wire [0:scan_right]      sov;

//64-bit core
//c64: if (regmode = 6) generate begin

/*
//table_start
?TABLE rom_instr LISTING(final) OPTIMIZE PARMS(ON-SET, OFF-SET);
*INPUTS*========*OUTPUTS*===============================================================================================*
|               |                                                                                                       |
| rom_addr_l2   | template                         ucode_end                                                            |
| |             | |                                | ucode_end_early                                                    |
| |             | |                                | | loop_begin                                                       |
| |             | |                                | | | loop_end                                                       |
| |             | |                                | | | | count_src                                                    | -- Can DC if not (loop_begin or loop_end)
| |             | |                                | | | | |                                                            |
| |             | |                                | | | | |    ext_rt                                                  |
| |             | |                                | | | | |    | ext_s1                                                |
| |             | |                                | | | | |    | | ext_s2                                              |
| |             | |                                | | | | |    | | | ext_s3                                            |
| |             | |                                | | | | |    | | | |                                                 |
| |             | |                                | | | | |    | | | |  sel0_5                                         |
| |             | |                                | | | | |    | | | |  | sel6_10                                      |
| |             | |                                | | | | |    | | | |  | |  sel11_15                                  |
| |             | |                                | | | | |    | | | |  | |  |  sel16_20                               |
| |             | |                                | | | | |    | | | |  | |  |  |  sel21_25                            |
| |             | |                                | | | | |    | | | |  | |  |  |  |  sel26_30                         |
| |             | |                                | | | | |    | | | |  | |  |  |  |  | sel31                          |
| |             | |                                | | | | |    | | | |  | |  |  |  |  | |                              |
| |             | |                                | | | | |    | | | |  | |  |  |  |  | |  cr_bf2fxm                   |
| |             | |                                | | | | |    | | | |  | |  |  |  |  | |  | skip_cond                 |
| |             | |                                | | | | |    | | | |  | |  |  |  |  | |  | | skip_zero               | -- Can DC if loop_begin not set
| |             | |                                | | | | |    | | | |  | |  |  |  |  | |  | | | skip_nop              | -- Optimize to only be in odd side
| |             | |                                | | | | |    | | | |  | |  |  |  |  | |  | | | | loop_addr           | -- Can DC if loop_end not set; always odd side
| |             | |                                | | | | |    | | | |  | |  |  |  |  | |  | | | | |          loop_init| -- 1 less than # of times to loop; Can DC if not loop_begin or not count_src=111
| |             | |                                | | | | |    | | | |  | |  |  |  |  | |  | | | | |          |   ep   |
| |             | |         1111111111222222222233 | | | | |    | | | |  | |  |  |  |  | |  | | | | |          |   |    |
| 0123456789    | 01234567890123456789012345678901 | | | | 012  | | | |  | 01 01 01 01 | |  | | | | 0123456789 012 |    |
*TYPE*==========+=======================================================================================================+
| PPPPPPPPPP    | SSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSS S S S S SSS  S S S S  S SS SS SS SS S S  S S S S SSSSSSSSSS SSS S    |
*OPTIMIZE*----->| AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA B B B B CCC  X X X X  X XX XX XX XX X X  X X X X XXXXXXXXXX XYX X    |
*TERMS*=========+=======================================================================================================+
| 0000000001    | 10001000001000000000000000000000 0 0 0 - ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # lbz s1,0(s0)
| 0000000011    | 01010000001000100100010000101110 0 0 0 - ---  1 1 1 -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # rlwimi s2,s1,8,16,23
| 0000000101    | 01111100010000100000101101111000 0 0 0 - ---  1 1 1 -  0 00 00 00 00 0 0  0 1 - 0 ---------- --- -    | # or s2,s2,s1 	-skip_c
| 0000000111    | 01101000000-----0000000000000000 1 - 0 - ---  0 1 - -  0 00 01 00 00 0 0  0 0 - 0 ---------- --- -    | # xori RA,s0,0

| 0000010001    | 01111100001-----000000001010111- 0 0 0 - ---  1 0 1 -  0 00 01 00 00 0 -  0 0 - 0 ---------- --- 1    | # lbzx s1,RA,s0
| 0000010011    | 01111100010-----000110001010111- 0 0 0 - ---  1 0 1 -  0 00 01 00 00 0 -  0 0 - 0 ---------- --- 1    | # lbzx s2,RA,s3
| 0000010101    | 01010100010000100100010000101110 0 0 0 - ---  1 1 - -  0 00 00 00 00 0 0  0 1 - 0 ---------- --- 0    | # rlwinm s2,s2,8,16,23 	-skip_c
| 0000010111    | 01101000010-----0000000000000000 0 1 0 - ---  0 1 - -  0 00 11 00 00 0 0  0 0 - 0 ---------- --- 0    | # xori RT,s2,0 	-end for non-update

| 0000100001    | 10001000001000000000000000000000 0 0 0 - ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # lbz s1,0(s0)
| 0000100011    | 01010000001000100100010000101110 0 0 0 - ---  1 1 1 -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # rlwimi s2,s1,8,16,23
| 0000100101    | 01111100010000100000101101111000 0 0 0 - ---  1 1 1 -  0 00 00 00 00 0 0  0 1 - 0 ---------- --- -    | # or s2,s2,s1 	-skip_c
| 0000100111    | 01101000000-----0000000000000000 1 - 0 - ---  0 1 - -  0 00 01 00 00 0 0  0 0 - 0 ---------- --- -    | # xori RA,s0,0

| 0000110001    | 0111110000000000-----01000010100 0 0 0 - ---  1 1 0 -  0 00 00 01 00 0 0  0 0 - 0 ---------- --- -    | # add s0,s0,RB
| 0000110011    | 10001000010000000000000000000001 0 0 0 - ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # lbz s2,1(s0)
| 0000110101    | 01010100010000100100010000101110 0 0 0 - ---  1 1 - -  0 00 00 00 00 0 0  0 1 - 0 ---------- --- -    | # rlwinm s2,s2,8,16,23 	-skip_c
| 0000110111    | 01111100010----------11100110100 0 1 0 - ---  0 1 - -  0 00 11 -- 00 0 0  0 0 - 0 ---------- --- -    | # extsh RT,s2 	-end for non-update

| 0001000001    | 10001000010000000000000000000000 0 0 0 - ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # lbz s2,0(s0)
| 0001000011    | 01010100010000100100000000111110 0 0 0 0 ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # rlwinm s2,s2,8,0,31
| 0001000101    | 01111100010000100000101101111000 0 0 0 1 111  1 1 1 -  0 00 00 00 00 0 0  0 0 - 0 0001000010 --- -    | # or s2,s2,s1 	-loop_end
| 0001000111    | 01010000010000101000010000101110 0 0 0 - ---  1 1 1 -  0 00 00 00 00 0 0  0 1 - 0 ---------- --- -    | # rlwimi s2,s2,16,16,23 	-skip_c
| 0001001001    | 01101000010-----0000000000000000 0 1 0 - ---  0 1 - -  0 00 11 00 00 0 0  0 0 - 0 ---------- --- -    | # xori RT,s2,0 	-end for non-update

| 0001010001    | 01111100010-----000000001010111- 0 0 0 - ---  1 0 1 -  0 00 01 00 00 0 -  0 0 - 0 ---------- --- 1    | # lbzx s2,RA,s0
| 0001010011    | 01010100010000100100000000111110 0 0 0 0 ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- 0    | # rlwinm s2,s2,8,0,31
| 0001010101    | 01111100010000100000101101111000 0 0 0 1 111  1 1 1 -  0 00 00 00 00 0 0  0 0 - 0 0001010010 --- 0    | # or s2,s2,s1 	-loop_end
| 0001010111    | 01010000010000101000010000101110 0 0 0 - ---  1 1 1 -  0 00 00 00 00 0 0  0 1 - 0 ---------- --- 0    | # rlwimi s2,s2,16,16,23 	-skip_c
| 0001011001    | 01101000010-----0000000000000000 0 1 0 - ---  0 1 - -  0 00 11 00 00 0 0  0 0 - 0 ---------- --- 0    | # xori RT,s2,0 	-end for non-update
| 0001011011    | 011111-----000010000001000010100 1 - 0 - ---  0 1 1 -  0 10 00 00 00 0 0  0 0 - 0 ---------- --- 0    | # add RA,s1,s0

| 0001100001    | 1000100001000000---------------- 0 - 0 - ---  1 1 - -  0 00 00 01 01 1 1  0 0 - 0 ---------- --- -    | # lbz s2,D(s0)
| 0001100011    | 01010100010000100100000000111110 0 - 0 0 ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # rlwinm s2,s2,8,0,31
| 0001100101    | 01111100010000100000101101111000 0 - 0 1 111  1 1 1 -  0 00 00 00 00 0 0  0 0 - 0 0001100010 --- -    | # or s2,s2,s1 	-loop_end
| 0001100111    | 01010000010000101000010000101110 0 - 0 - ---  1 1 1 -  0 00 00 00 00 0 0  0 1 - 0 ---------- --- -    | # rlwimi s2,s2,16,16,23 	-skip_c
| 0001101001    | 01111100010----------11110110100 1 - 0 - ---  0 1 - -  0 00 11 -- 00 0 0  0 0 - 0 ---------- --- -    | # extsw RT,s2

| 0001110001    | 01111100010-----000000001010111- 0 0 0 - ---  1 0 1 -  0 00 01 00 00 0 -  0 0 - 0 ---------- --- -    | # lbzx s2,RA,s0
| 0001110011    | 01010100010000100100000000111110 0 0 0 0 ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # rlwinm s2,s2,8,0,31
| 0001110101    | 01111100010000100000101101111000 0 0 0 1 111  1 1 1 -  0 00 00 00 00 0 0  0 0 - 0 0001110010 --- -    | # or s2,s2,s1 	-loop_end
| 0001110111    | 01010000010000101000010000101110 0 0 0 - ---  1 1 1 -  0 00 00 00 00 0 0  0 1 - 0 ---------- --- -    | # rlwimi s2,s2,16,16,23 	-skip_c
| 0001111001    | 01111100010----------11110110100 0 1 0 - ---  0 1 - -  0 00 11 -- 00 0 0  0 0 - 0 ---------- --- -    | # extsw RT,s2 	-end for non-update
| 0001111011    | 011111-----000010000001000010100 1 - 0 - ---  0 1 1 -  0 10 00 00 00 0 0  0 0 - 0 ---------- --- -    | # add RA,s1,s0

| 0010000001    | 10001000010000000000000000000000 0 0 0 - ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # lbz s2,0(s0)
| 0010000011    | 01111000010000100100010111100100 0 0 0 0 ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # rldicr s2,s2,8,55
| 0010000101    | 01111100010000100000101101111000 0 0 0 1 111  1 1 1 -  0 00 00 00 00 0 0  0 0 - 0 0010000010 --- -    | # or s2,s2,s1 	-loop_end
| 0010000111    | 01111000001000010100000000000000 0 0 0 0 ---  1 1 - -  0 00 00 00 00 0 0  0 1 - 0 ---------- --- -    | # rldicl s1,s1,8,0 	-skip_c
| 0010001001    | 00111000010000010000000000000000 0 0 0 - 111  1 1 - -  0 00 00 00 00 0 0  0 1 - 0 0010000110 --- -    | # addi s2,s1,0 	-skip_c
| 0010001011    | 001110-------------------------0 1 - 0 - ---  0 0 - -  0 10 01 01 01 1 0  0 0 - 0 ---------- --- -    | # addi RA,RA,DS

| 0010010001    | 01111100010-----000000001010111- 0 0 0 - ---  1 0 1 -  0 00 01 00 00 0 -  0 0 - 0 ---------- --- 1    | # lbzx s2,RA,s0
| 0010010011    | 01111000010000100100010111100100 0 0 0 0 ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- 0    | # rldicr s2,s2,8,55
| 0010010101    | 01111100010000100000101101111000 0 0 0 1 111  1 1 1 -  0 00 00 00 00 0 0  0 0 - 0 0010010010 --- 0    | # or s2,s2,s1 	-loop_end
| 0010010111    | 01111000001000010100000000000000 0 0 0 0 ---  1 1 - -  0 00 00 00 00 0 0  0 1 - 0 ---------- --- 0    | # rldicl s1,s1,8,0 	-skip_c
| 0010011001    | 00111000010000010000000000000000 0 0 0 - 111  1 1 - -  0 00 00 00 00 0 0  0 1 - 0 0010010110 --- 0    | # addi s2,s1,0 	-skip_c
| 0010011011    | 00111000001-----1111111111111001 0 - 0 - ---  1 0 - -  0 00 01 00 00 0 0  0 0 - 0 ---------- --- 0    | # addi s1,RA,-7

| 0010100001    | -------------------------------- 0 - 0 - ---  - - - -  - -- -- -- -- - -  0 - - 1 ---------- --- -    | # nop
| 0010100011    | 00111000000000000000000000000100 0 - 0 1 100  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 0010100010 --- -    | # addi s0,s0,4 	-loop_end

| 0010110001    | -------------------------------- 0 - 0 - ---  - - - -  - -- -- -- -- - -  0 - - 1 ---------- --- -    | # nop
| 0010110011    | 01010100010000101100000000111110 0 - 0 0 ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # rlwinm s2,s2,24,0,31
| 0010110101    | 01010000001000101000001000011110 0 - 0 0 ---  1 1 1 -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # rlwimi s2,s1,16,8,15
| 0010110111    | 01010000001000100100010000101110 0 - 0 0 ---  1 1 1 -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # rlwimi s2,s1,8,16,23
| 0010111001    | 00111000000000000000000000000100 0 - 0 0 ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # addi s0,s0,4
| 0010111011    | -------------------------------- 0 - 0 - 101  - - - -  - -- -- -- -- - -  0 - - 1 0010110010 --- -    | # nop
| 0010111101    | 01010100010000100100000000101110 0 - 0 0 ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # rlwinm s2,s2,8,0,23
| 0010111111    | 01111100010000100000101101111000 0 - 0 1 000  1 1 1 -  0 00 00 00 00 0 0  0 0 - 0 0010111100 --- -    | # or s2,s2,s1 	-loop_end
| 0011000001    | -------------------------------- 0 - 0 1 001  - - - -  - -- -- -- -- - -  0 - - 1 0011000000 --- -    | # nop         -loop_end

| 0011010001    | 00111000000-----0000000000000000 0 - 0 - ---  1 0 - -  0 00 01 00 00 0 0  0 0 - 0 ---------- --- -    | # addi s0,RA,0
| 0011010011    | 00111000000000000000000000000001 0 - 0 0 ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # addi s0,s0,1
| 0011010101    | 0111110000100000-----0001010111- 0 - 0 0 ---  1 1 0 -  0 00 00 01 00 0 -  0 0 - 0 ---------- --- -    | # lbzx s1,s0,RB
| 0011010111    | 01010000001000101000001000011110 0 - 0 0 ---  1 1 1 -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # rlwimi s2,s1,16,8,15
| 0011011001    | 00111000000000000000000000000001 0 - 0 0 ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # addi s0,s0,1
| 0011011011    | 0111110000100000-----0001010111- 0 - 0 0 ---  1 1 0 -  0 00 00 01 00 0 -  0 0 - 0 ---------- --- -    | # lbzx s1,s0,RB
| 0011011101    | 01111100010-----0000101101111000 0 - 0 1 110  0 1 1 -  0 00 11 00 00 0 0  0 0 - 0 0011010010 --- -    | # or RT,s2,s1 	-loop_end
| 0011011111    | 01010100010000100100000000101110 0 - 0 0 ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # rlwinm s2,s2,8,0,23
| 0011100001    | 01111100010000100000101101111000 0 - 0 1 010  1 1 1 -  0 00 00 00 00 0 0  0 0 - 0 0011011110 --- -    | # or s2,s2,s1 	-loop_end
| 0011100011    | -------------------------------- 0 - 0 1 011  - - - -  - -- -- -- -- - -  0 - - 1 0011100010 --- -    | # nop         -loop_end


| 0100000001    | 00111000000--------------------- 0 0 0 - ---  1 0 - -  0 00 01 01 01 1 1  0 0 - 0 ---------- --- -    | # addi s0,RA,D
| 0100000011    | 010100-----000100000011000111110 0 0 0 - ---  1 0 1 -  0 01 00 00 00 0 0  0 1 - 0 ---------- --- -    | # rlwimi s2,RS,0,24,31 	-skip_c
| 0100000101    | 01010100010000100100000000111110 0 0 0 - ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # rlwinm s2,s2,8,0,31
| 0100000111    | 001110-------------------------- 1 - 0 - ---  0 0 - -  0 10 01 01 01 1 1  0 0 - 0 ---------- --- -    | # addi RA,RA,D

| 0100010001    | 00111000000-----0000000000000001 0 0 0 - ---  1 0 - -  0 00 01 00 00 0 0  0 0 - 0 ---------- --- 0    | # addi s0,RA,1
| 0100010011    | 010100-----000100000011000111110 0 0 0 - ---  1 0 1 -  0 01 00 00 00 0 0  0 1 - 0 ---------- --- 0    | # rlwimi s2,RS,0,24,31 	-skip_c
| 0100010101    | 01010100010000100100000000111110 0 0 0 - ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- 0    | # rlwinm s2,s2,8,0,31
| 0100010111    | 00111000000-----0000000000000000 0 - 0 - ---  1 0 - -  0 00 01 00 00 0 0  0 0 - 0 ---------- --- 0    | # addi s0,RA,0

| 0101000001    | 010101-----000100000000000111110 0 0 0 - ---  1 0 - -  0 01 00 00 00 0 0  0 1 - 0 ---------- --- -    | # rlwinm s2,RS,0,0,31 	-skip_c
| 0101000011    | 010100-----000101000000000001110 0 0 0 - ---  1 0 1 -  0 01 00 00 00 0 0  0 1 - 0 ---------- --- -    | # rlwimi s2,RS,16,0,7 	-skip_c
| 0101000101    | 10011000010000000000000000000000 0 0 0 - ---  - 1 - 1  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # stb s2,0(s0)
| 0101000111    | 01010100010000100100000000111110 0 0 0 0 ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # rlwinm s2,s2,8,0,31
| 0101001001    | 001110-------------------------- 1 - 0 - 111  0 0 - -  0 10 01 01 01 1 1  0 0 - 0 0101000110 --- -    | # addi RA,RA,D

| 0101010001    | 010101-----000100000000000111110 0 0 0 - ---  1 0 - -  0 01 00 00 00 0 0  0 1 - 0 ---------- --- 0    | # rlwinm s2,RS,0,0,31 	-skip_c
| 0101010011    | 010100-----000101000000000001110 0 0 0 - ---  1 0 1 -  0 01 00 00 00 0 0  0 1 - 0 ---------- --- 0    | # rlwimi s2,RS,16,0,7 	-skip_c
| 0101010101    | 0111110001000000-----0011010111- 0 0 0 - ---  - 1 0 1  0 00 00 01 00 0 -  0 0 - 0 ---------- --- 1    | # stbx s2,s0,RB
| 0101010111    | 01010100010000100100000000111110 0 0 0 0 ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- 0    | # rlwinm s2,s2,8,0,31
| 0101011001    | 011111---------------01000010100 1 - 0 - 111  0 0 0 -  0 10 01 01 00 0 0  0 0 - 0 0101010110 --- 0    | # add RA,RA,RB

| 0110000001    | 00111000000-----0000000000000000 0 0 0 - ---  1 0 - -  0 00 01 00 00 0 0  0 0 - 0 ---------- --- -    | # addi s0,RA,0
| 0110000011    | 01111000001000010100000000000000 0 0 0 0 ---  1 1 - -  0 00 00 00 00 0 0  0 1 - 0 ---------- --- -    | # rldicl s1,s1,8,0 	-skip_c
| 0110000101    | 01111000001000100100000000000000 0 0 0 - 111  1 1 - -  0 00 00 00 00 0 0  0 1 - 0 0110000010 --- -    | # rldicl s2,s1,8,0 	-skip_c
| 0110000111    | 00111000000000000000000000000001 0 0 0 0 ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # addi s0,s0,1
| 0110001001    | 1001100001000000---------------0 0 1 0 - 111  - 1 - 1  0 00 00 01 01 1 0  0 0 - 0 0110000110 --- -    | # stb s2,DS(s0) 	-end for non-update

| 0110010001    | 00111000000-----0000000000000000 0 0 0 - ---  1 0 - -  0 00 01 00 00 0 0  0 0 - 0 ---------- --- 0    | # addi s0,RA,0
| 0110010011    | 01111000001000010100000000000000 0 0 0 0 ---  1 1 - -  0 00 00 00 00 0 0  0 1 - 0 ---------- --- 0    | # rldicl s1,s1,8,0 	-skip_c
| 0110010101    | 01111000001000100100000000000000 0 0 0 - 111  1 1 - -  0 00 00 00 00 0 0  0 1 - 0 0110010010 --- 0    | # rldicl s2,s1,8,0 	-skip_c
| 0110010111    | 00111000000000000000000000000001 0 0 0 0 ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- 0    | # addi s0,s0,1
| 0110011001    | 0111110001000000-----0011010111- 0 1 0 - 111  - 1 0 1  0 00 00 01 00 0 -  0 0 - 0 0110010110 --- 1    | # stbx s2,s0,RB 	-end for non-update


| 0110100001    | -------------------------------- 0 - 0 - ---  - - - -  - -- -- -- -- - -  0 - - 1 ---------- --- -    | # nop
| 0110100011    | 00111000000000000000000000000100 0 - 0 1 100  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 0110100010 --- -    | # addi s0,s0,4 	-loop_end

| 0110110001    | -------------------------------- 0 - 0 - ---  - - - -  - -- -- -- -- - -  0 - - 1 ---------- --- -    | # nop
| 0110110011    | 10011000010000000000000000000000 0 - 0 0 ---  - 1 - 1  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # stb s2,0(s0)
| 0110110101    | 10011000010000000000000000000001 0 - 0 0 ---  - 1 - 1  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # stb s2,1(s0)
| 0110110111    | 10011000010000000000000000000010 0 - 0 0 ---  - 1 - 1  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # stb s2,2(s0)
| 0110111001    | 10011000010000000000000000000011 0 - 0 0 ---  - 1 - 1  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # stb s2,3(s0)
| 0110111011    | -------------------------------- 0 - 0 - 101  - - - -  - -- -- -- -- - -  0 - - 1 0110110010 --- -    | # nop
| 0110111101    | -------------------------------- 0 - 0 - ---  - - - -  - -- -- -- -- - -  0 - - 1 ---------- --- -    | # nop
| 0110111111    | 00111000000000000000000000000001 0 - 0 0 ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # addi s0,s0,1
| 0111000001    | -------------------------------- - - 0 - 000  - - - -  - -- -- -- -- - -  0 - - - 0110111110 --- -    | # nop

| 0111010001    | -------------------------------- 0 - 0 - ---  - - - -  - -- -- -- -- - -  0 - - 1 ---------- --- -    | # nop
| 0111010011    | 0111110001000000-----0011010111- 0 - 0 0 ---  - 1 0 1  0 00 00 01 00 0 -  0 0 - 0 ---------- --- -    | # stbx s2,s0,RB
| 0111010101    | 01010100010000100100000000111110 0 - 0 0 ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # rlwinm s2,s2,8,0,31
| 0111010111    | 00111000000000000000000000000001 0 - 0 0 ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # addi s0,s0,1
| 0111011001    | 0111110001000000-----0011010111- 0 - 0 0 ---  - 1 0 1  0 00 00 01 00 0 -  0 0 - 0 ---------- --- -    | # stbx s2,s0,RB
| 0111011011    | 01010100010000100100000000111110 0 - 0 0 ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # rlwinm s2,s2,8,0,31
| 0111011101    | 00111000000000000000000000000001 0 - 0 1 110  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 0111010010 --- -    | # addi s0,s0,1 	-loop_end
| 0111011111    | -------------------------------- 0 - 0 - ---  - - - -  - -- -- -- -- - -  0 - - 1 ---------- --- -    | # nop
| 0111100001    | 00111000000000000000000000000001 0 - 0 0 ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # addi s0,s0,1
| 0111100011    | 01100000000000000000000000000000 1 - 0 - 010  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 0111100000 --- -    | # ori 0,0,0 (nop)


| 0101100001    | 01010100000000010000000000000110 0 - 0 - ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # rlwinm s1,s0,0,0,3
| 0101100011    | 01010100001000001110000100111110 0 - 0 - ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # srwi s0,s1,4
| 0101100101    | 01010100001000001100001000111110 0 - 0 - ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # srwi s0,s1,8
| 0101100111    | 01010100001000001000010000111110 0 - 0 - ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # srwi s0,s1,16
| 0101101001    | 01111100001----------0010010000- 0 - 0 - ---  - 1 - -  0 00 01 01 00 0 -  1 0 - 0 ---------- --- -    | # mtocrf BF,s1

| 0101110001    | 01111100000101000000-0000010011- 0 - 0 - ---  1 - - -  0 00 00 00 00 0 -  0 0 - 0 ---------- --- -    | # mfocrf s0,0x40
| 0101110011    | 01111100000100100000-0000010011- 0 - 0 - ---  1 - - -  0 00 00 00 00 0 -  0 0 - 0 ---------- --- -    | # mfocrf s0,0x20
| 0101110101    | 01111100000100010000-0000010011- 0 - 0 - ---  1 - - -  0 00 00 00 00 0 -  0 0 - 0 ---------- --- -    | # mfocrf s0,0x10
| 0101110111    | 01111100000100001000-0000010011- 0 - 0 - ---  1 - - -  0 00 00 00 00 0 -  0 0 - 0 ---------- --- -    | # mfocrf s0,0x08
| 0101111001    | 01111100000100000100-0000010011- 0 - 0 - ---  1 - - -  0 00 00 00 00 0 -  0 0 - 0 ---------- --- -    | # mfocrf s0,0x04
| 0101111011    | 01111100000100000010-0000010011- 0 - 0 - ---  1 - - -  0 00 00 00 00 0 -  0 0 - 0 ---------- --- -    | # mfocrf s0,0x02
| 0101111101    | 01111100000100000001-0000010011- 0 - 0 - ---  1 - - -  0 00 00 00 00 0 -  0 0 - 0 ---------- --- -    | # mfocrf s0,0x01


| 0111110001    | 011111-----101000000-0010010000- 0 - 0 - ---  - 0 - -  0 01 00 00 00 0 -  0 0 - 0 ---------- --- -    | # mtocrf 0x40,RS
| 0111110011    | 011111-----100010000-0010010000- 0 - 0 - ---  - 0 - -  0 01 00 00 00 0 -  0 0 - 0 ---------- --- -    | # mtocrf 0x10,RS
| 0111110101    | 011111-----100000100-0010010000- 0 - 0 - ---  - 0 - -  0 01 00 00 00 0 -  0 0 - 0 ---------- --- -    | # mtocrf 0x04,RS
| 0111110111    | 011111-----100000001-0010010000- 1 - 0 - ---  - 0 - -  0 01 00 00 00 0 -  0 0 - 0 ---------- --- -    | # mtocrf 0x01,RS



| 1010100001    | 001110-------------------------- 1 - 0 - ---  0 0 - -  0 10 01 01 01 1 1  0 0 - 0 ---------- --- -    | # addi RA,RA,D

| 1010101001    | 100010-----000000000000000000000 0 - 0 - ---  0 1 - -  0 01 00 00 00 0 0  0 0 - 0 ---------- --- -    | # lbz RT,0(s0)

| 1010110001    | 001110-------------------------- 1 - 0 - ---  0 0 - -  0 10 01 01 01 1 1  0 0 - 0 ---------- --- -    | # addi RA,RA,D

| 1010111001    | 101000-----000000000000000000000 0 - 0 - ---  0 1 - -  0 01 00 00 00 0 0  0 0 - 0 ---------- --- -    | # lhz RT,0(s0)

| 1011000001    | 001110-------------------------- 1 - 0 - ---  0 0 - -  0 10 01 01 01 1 1  0 0 - 0 ---------- --- -    | # addi RA,RA,D

| 1011001001    | 100000-----000000000000000000000 0 - 0 - ---  0 1 - -  0 01 00 00 00 0 0  0 0 - 0 ---------- --- -    | # lwz RT,0(s0)

| 1011010001    | 001110-------------------------0 1 - 0 - ---  0 0 - -  0 10 01 01 01 1 0  0 0 - 0 ---------- --- -    | # addi RA,RA,DS

| 1011011001    | 111010-----000000000000000000000 0 - 0 - ---  0 1 - -  0 01 00 00 00 0 0  0 0 - 0 ---------- --- -    | # ld RT,0(s0)

| 1011100001    | 001110-------------------------- 1 - 0 - ---  0 0 - -  0 10 01 01 01 1 1  0 0 - 0 ---------- --- -    | # addi RA,RA,D

| 1011101001    | 101010-----000000000000000000000 0 - 0 - ---  0 1 - -  0 01 00 00 00 0 0  0 0 - 0 ---------- --- -    | # lha RT,0(s0)

| 1011111001    | 111010-----000000000000000000010 0 - 0 - ---  0 1 - -  0 01 00 00 00 0 0  0 0 - 0 ---------- --- -    | # lwa RT,0(s0)



| 1000110001    | 01111100010-----000000001010111- 0 - 0 - ---  1 0 1 -  0 00 01 00 00 0 -  0 0 - 0 ---------- --- -    | # lbzx s2,RA,s0
| 1000110011    | 01010100010000100100000000111110 0 - 0 0 ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # rlwinm s2,s2,8,0,31
| 1000110101    | 01111100010000100000101101111000 0 - 0 1 111  1 1 1 -  0 00 00 00 00 0 0  0 0 - 0 1000110010 --- -    | # or s2,s2,s1 	-loop_end
| 1000110111    | 01010000010000101000010000101110 0 - 0 - ---  1 1 1 -  0 00 00 00 00 0 0  0 1 - 0 ---------- --- -    | # rlwimi s2,s2,16,16,23 	-skip_c
| 1000111001    | 011111-----000000001010011111000 1 - 0 - ---  0 - 1 -  0 01 00 00 00 0 0  0 0 - 0 ---------- --- -    | # mfifgpr RT,s2,0 	-end

| 1001110001    | 01111100010-----000000001010111- 0 - 0 - ---  1 0 1 -  0 00 01 00 00 0 -  0 0 - 0 ---------- --- -    | # lbzx s2,RA,s0
| 1001110011    | 01010100010000100100000000111110 0 - 0 0 ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # rlwinm s2,s2,8,0,31
| 1001110101    | 01111100010000100000101101111000 0 - 0 1 111  1 1 1 -  0 00 00 00 00 0 0  0 0 - 0 1001110010 --- -    | # or s2,s2,s1 	-loop_end
| 1001110111    | 01010000010000101000010000101110 0 - 0 - ---  1 1 1 -  0 00 00 00 00 0 0  0 1 - 0 ---------- --- -    | # rlwimi s2,s2,16,16,23 	-skip_c
| 1001111001    | 011111-----000000001010011111010 1 - 0 - ---  0 - 1 -  0 01 00 00 00 0 0  0 0 - 0 ---------- --- -    | # mfixfgpr RT,s2,0 	-end

| 1001000001    | 10001000010000000000000000000000 0 0 0 - ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # lbz s2,0(s0)
| 1001000011    | 01010100010000100100000000111110 0 0 0 0 ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # rlwinm s2,s2,8,0,31
| 1001000101    | 01111100010000100000101101111000 0 0 0 1 111  1 1 1 -  0 00 00 00 00 0 0  0 0 - 0 1001000010 --- -    | # or s2,s2,s1 	-loop_end
| 1001000111    | 01010000010000101000010000101110 0 0 0 - ---  1 1 1 -  0 00 00 00 00 0 0  0 1 - 0 ---------- --- -    | # rlwimi s2,s2,16,16,23 	-skip_c
| 1001001001    | 01111100000000000001010011111100 0 1 0 - ---  0 - 1 -  0 01 00 00 00 0 0  0 0 - 0 ---------- --- -    | # mfsfgpr RT,s2,0 	-end for non-update

| 1001010001    | 01111100010-----000000001010111- 0 0 0 - ---  1 0 1 -  0 00 01 00 00 0 -  0 0 - 0 ---------- --- -    | # lbzx s2,RA,s0
| 1001010011    | 01010100010000100100000000111110 0 0 0 0 ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # rlwinm s2,s2,8,0,31
| 1001010101    | 01111100010000100000101101111000 0 0 0 1 111  1 1 1 -  0 00 00 00 00 0 0  0 0 - 0 1001010010 --- -    | # or s2,s2,s1 	-loop_end
| 1001010111    | 01010000010000101000010000101110 0 0 0 - ---  1 1 1 -  0 00 00 00 00 0 0  0 1 - 0 ---------- --- -    | # rlwimi s2,s2,16,16,23 	-skip_c
| 1001011001    | 011111-----000000001010011111100 0 1 0 - ---  0 - 1 -  0 01 00 00 00 0 0  0 0 - 0 ---------- --- -    | # mfsfgpr RT,s2,0 	-end for non-update
| 1001011011    | 011111-----000010000001000010100 1 - 0 - ---  0 1 1 -  0 10 00 00 00 0 0  0 0 - 0 ---------- --- -    | # add RA,s1,s0

| 1010000001    | 10001000010000000000000000000000 0 0 0 - ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # lbz s2,0(s0)
| 1010000011    | 01111000010000100100010111100100 0 0 0 0 ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # rldicr s2,s2,8,55
| 1010000101    | 01111100010000100000101101111000 0 0 0 1 111  1 1 1 -  0 00 00 00 00 0 0  0 0 - 0 1010000010 --- -    | # or s2,s2,s1 	-loop_end
| 1010000111    | 01111000001000010100000000000000 0 0 0 0 ---  1 1 - -  0 00 00 00 00 0 0  0 1 - 0 ---------- --- -    | # rldicl s1,s1,8,0 	-skip_c
| 1010001001    | 01101000001000100000000000000000 0 0 0 - 111  1 1 - -  0 00 00 00 00 0 0  0 1 - 0 1010000110 --- -    | # xori s2,s1,0 	-skip_c
| 1010001011    | 001110-------------------------- 1 - 0 - ---  0 0 - -  0 10 01 01 01 1 1  0 0 - 0 ---------- --- -    | # addi RA,RA,D

| 1010010001    | 01111100010-----000000001010111- 0 0 0 - ---  1 0 1 -  0 00 01 00 00 0 -  0 0 - 0 ---------- --- 1    | # lbzx s2,RA,s0
| 1010010011    | 01111000010000100100010111100100 0 0 0 0 ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- 0    | # rldicr s2,s2,8,55
| 1010010101    | 01111100010000100000101101111000 0 0 0 1 111  1 1 1 -  0 00 00 00 00 0 0  0 0 - 0 1010010010 --- 0    | # or s2,s2,s1 	-loop_end
| 1010010111    | 01111000001000010100000000000000 0 0 0 0 ---  1 1 - -  0 00 00 00 00 0 0  0 1 - 0 ---------- --- 0    | # rldicl s1,s1,8,0 	-skip_c
| 1010011001    | 01101000001000100000000000000000 0 0 0 - 111  1 1 - -  0 00 00 00 00 0 0  0 1 - 0 1010010110 --- 0    | # xori s2,s1,0 	-skip_c
| 1010011011    | 00111000001-----1111111111111001 0 - 0 - ---  1 0 - -  0 00 01 00 00 0 0  0 0 - 0 ---------- --- 0    | # addi s1,RA,-7

| 1100110001    | 00111000000-----0000000000000000 0 - 0 - ---  1 0 - -  0 00 01 00 00 0 0  0 0 - 0 ---------- --- -    | # addi s0,RA,0
| 1100110011    | 01010100001000100000000000111110 0 - 0 - ---  1 1 - -  0 00 00 00 00 0 0  0 1 - 0 ---------- --- -    | # rlwinm s2,s1,0,0,31 	-skip_c
| 1100110101    | 01010000001000101000000000001110 0 - 0 - ---  1 1 1 -  0 00 00 00 00 0 0  0 1 - 0 ---------- --- -    | # rlwimi s2,s1,16,0,7 	-skip_c
| 1100110111    | 00111000000000000000000000000001 0 - 0 0 ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # addi s0,s0,1
| 1100111001    | 0111110001000000-----0011010111- 1 - 0 - 111  - 1 0 1  0 00 00 01 00 0 -  0 0 - 0 1100110110 --- -    | # stbx s2,s0,RB

| 1101000001    | 00111000000--------------------- 0 0 0 - ---  1 0 - -  0 00 01 01 01 1 1  0 0 - 0 ---------- --- -    | # addi s0,RA,D
| 1101000011    | 01010100001000100000000000111110 0 0 0 - ---  1 1 - -  0 00 00 00 00 0 0  0 1 - 0 ---------- --- -    | # rlwinm s2,s1,0,0,31 	-skip_c
| 1101000101    | 01010000001000101000000000001110 0 0 0 - ---  1 1 1 -  0 00 00 00 00 0 0  0 1 - 0 ---------- --- -    | # rlwimi s2,s1,16,0,7 	-skip_c
| 1101000111    | 00111000000000000000000000000001 0 0 0 0 ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # addi s0,s0,1
| 1101001001    | 10011000010000000000000000000000 0 1 0 - 111  - 1 - 1  0 00 00 00 00 0 0  0 0 - 0 1101000110 --- -    | # stb s2,0(s0) 	-end for non-update

| 1101010001    | 00111000000-----0000000000000000 0 0 0 - ---  1 0 - -  0 00 01 00 00 0 0  0 0 - 0 ---------- --- -    | # addi s0,RA,0
| 1101010011    | 01010100001000100000000000111110 0 0 0 - ---  1 1 - -  0 00 00 00 00 0 0  0 1 - 0 ---------- --- -    | # rlwinm s2,s1,0,0,31 	-skip_c
| 1101010101    | 01010000001000101000000000001110 0 0 0 - ---  1 1 1 -  0 00 00 00 00 0 0  0 1 - 0 ---------- --- -    | # rlwimi s2,s1,16,0,7 	-skip_c
| 1101010111    | 00111000000000000000000000000001 0 0 0 0 ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # addi s0,s0,1
| 1101011001    | 0111110001000000-----0011010111- 0 1 0 - 111  - 1 0 1  0 00 00 01 00 0 -  0 0 - 0 1101010110 --- -    | # stbx s2,s0,RB 	-end for non-update

| 1110000001    | 01111000001000100100000000000000 0 0 0 - ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # rldicl s2,s1,8,0
| 1110000011    | 01111000001000010100000000000000 0 0 0 0 ---  1 1 - -  0 00 00 00 00 0 0  0 1 - 0 ---------- --- -    | # rldicl s1,s1,8,0 	-skip_c
| 1110000101    | 01111000001000100100000000000000 0 0 0 - 111  1 1 - -  0 00 00 00 00 0 0  0 1 - 0 1110000010 --- -    | # rldicl s2,s1,8,0 	-skip_c
| 1110000111    | 1001100001000000---------------- 0 0 0 - ---  - 1 - 1  0 00 00 01 01 1 1  0 0 - 0 ---------- --- -    | # stb s2,D(s0)
| 1110001001    | 01111000010000100100000000000000 0 0 0 0 ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # rldicl s2,s2,8,0
| 1110001011    | 001110-------------------------- 1 - 0 - 111  0 0 - -  0 10 01 01 01 1 1  0 0 - 0 1110001000 --- -    | # addi RA,RA,D

| 1110010001    | 01111000001000100100000000000000 0 0 0 - ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- 0    | # rldicl s2,s1,8,0
| 1110010011    | 01111000001000010100000000000000 0 0 0 0 ---  1 1 - -  0 00 00 00 00 0 0  0 1 - 0 ---------- --- 0    | # rldicl s1,s1,8,0 	-skip_c
| 1110010101    | 01111000001000100100000000000000 0 0 0 - 111  1 1 - -  0 00 00 00 00 0 0  0 1 - 0 1110010010 --- 0    | # rldicl s2,s1,8,0 	-skip_c
| 1110010111    | 0111110001000000-----0011010111- 0 0 0 - ---  - 1 0 1  0 00 00 01 00 0 -  0 0 - 0 ---------- --- 1    | # stbx s2,s0,RB
| 1110011001    | 01111000010000100100000000000000 0 0 0 0 ---  1 1 - -  0 00 00 00 00 0 0  0 0 - 0 ---------- --- 0    | # rldicl s2,s2,8,0
| 1110011011    | 011111---------------01000010100 1 - 0 - 111  0 0 0 -  0 10 01 01 00 0 0  0 0 - 0 1110011000 --- 0    | # add RA,RA,RB



| 1111000001    | 001110-------------------------- 1 - 0 - ---  0 0 - -  0 10 01 01 01 1 1  0 0 - 0 ---------- --- -    | # addi RA,RA,DS

| 1111001001    | 110000-----000000000000000000000 0 - 0 - ---  0 1 - -  0 01 00 00 00 0 0  0 0 - 0 ---------- --- -    | # lfs FRT,0(s0)

| 1111010001    | 001110-------------------------- 1 - 0 - ---  0 0 - -  0 10 01 01 01 1 1  0 0 - 0 ---------- --- -    | # addi RA,RA,DS

| 1111011001    | 110010-----000000000000000000000 0 - 0 - ---  0 1 - -  0 01 00 00 00 0 0  0 0 - 0 ---------- --- -    | # lfd FRT,0(s0)


| 1100000001    | ----------------00001----------- 1 - 0 - ---  0 0 1 0  1 01 01 00 01 1 1  0 0 - 0 ---------- --- -    | # vvvvv FT,FA,FC,s1    - Original qpx op except B

| 1100001001    | 11111100010---------------100000 0 - 0 - ---  1 0 0 0  0 00 -- 11 -- 0 0  0 0 - 0 ---------- --- -    | # prenrm s2,FA         - prenorm both DP, SP

| 1100010001    | ----------------00001----------- 1 - 0 - ---  0 0 1 0  1 01 01 00 01 1 1  0 0 - 0 ---------- --- -    | # vvvvv FT,FA,FC,s1    - Original qpx op except B
*END*===========+=======================================================================================================+
?TABLE END rom_instr;
//table_end
*/

//assign_start

assign rom_instr_pt[1] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] ,
    rom_addr_l2[3] , rom_addr_l2[4] ,
    rom_addr_l2[5] , rom_addr_l2[6] ,
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 8'b01000000);
assign rom_instr_pt[2] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] ,
    rom_addr_l2[3] , rom_addr_l2[4] ,
    rom_addr_l2[5] , rom_addr_l2[6] ,
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 8'b00110000);
assign rom_instr_pt[3] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] ,
    rom_addr_l2[4] , rom_addr_l2[5] ,
    rom_addr_l2[6] , rom_addr_l2[7] ,
    rom_addr_l2[8] }) === 7'b1010000);
assign rom_instr_pt[4] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] ,
    rom_addr_l2[3] , rom_addr_l2[5] ,
    rom_addr_l2[6] , rom_addr_l2[7] ,
    rom_addr_l2[8] }) === 7'b0010000);
assign rom_instr_pt[5] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[3] , rom_addr_l2[5] ,
    rom_addr_l2[6] , rom_addr_l2[7] ,
    rom_addr_l2[8] }) === 7'b1110000);
assign rom_instr_pt[6] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] ,
    rom_addr_l2[3] , rom_addr_l2[4] ,
    rom_addr_l2[5] , rom_addr_l2[6] ,
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 8'b01001000);
assign rom_instr_pt[7] =
    (({ rom_addr_l2[1] , rom_addr_l2[4] ,
    rom_addr_l2[5] , rom_addr_l2[6] ,
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 6'b001000);
assign rom_instr_pt[8] =
    (({ rom_addr_l2[2] , rom_addr_l2[4] ,
    rom_addr_l2[5] , rom_addr_l2[6] ,
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 6'b111000);
assign rom_instr_pt[9] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[4] , rom_addr_l2[5] ,
    rom_addr_l2[6] , rom_addr_l2[7] ,
    rom_addr_l2[8] }) === 7'b0111000);
assign rom_instr_pt[10] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] ,
    rom_addr_l2[3] , rom_addr_l2[5] ,
    rom_addr_l2[6] , rom_addr_l2[7] ,
    rom_addr_l2[8] }) === 7'b0011000);
assign rom_instr_pt[11] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[3] , rom_addr_l2[5] ,
    rom_addr_l2[6] , rom_addr_l2[7] ,
    rom_addr_l2[8] }) === 7'b0011000);
assign rom_instr_pt[12] =
    (({ rom_addr_l2[0] , rom_addr_l2[2] ,
    rom_addr_l2[5] , rom_addr_l2[6] ,
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 6'b101000);
assign rom_instr_pt[13] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[2] , rom_addr_l2[3] ,
    rom_addr_l2[4] , rom_addr_l2[6] ,
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 8'b01110000);
assign rom_instr_pt[14] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[3] , rom_addr_l2[4] ,
    rom_addr_l2[6] , rom_addr_l2[7] ,
    rom_addr_l2[8] }) === 7'b0110000);
assign rom_instr_pt[15] =
    (({ rom_addr_l2[0] , rom_addr_l2[2] ,
    rom_addr_l2[3] , rom_addr_l2[4] ,
    rom_addr_l2[6] , rom_addr_l2[7] ,
    rom_addr_l2[8] }) === 7'b0101000);
assign rom_instr_pt[16] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[2] , rom_addr_l2[4] ,
    rom_addr_l2[6] , rom_addr_l2[7] ,
    rom_addr_l2[8] }) === 7'b0011000);
assign rom_instr_pt[17] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[2] , rom_addr_l2[3] ,
    rom_addr_l2[6] , rom_addr_l2[7] ,
    rom_addr_l2[8] }) === 7'b1000000);
assign rom_instr_pt[18] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[3] , rom_addr_l2[6] ,
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 6'b010000);
assign rom_instr_pt[19] =
    (({ rom_addr_l2[1] , rom_addr_l2[3] ,
    rom_addr_l2[6] , rom_addr_l2[7] ,
    rom_addr_l2[8] }) === 5'b10000);
assign rom_instr_pt[20] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] ,
    rom_addr_l2[3] , rom_addr_l2[6] ,
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 6'b111000);
assign rom_instr_pt[21] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[6] , rom_addr_l2[7] ,
    rom_addr_l2[8] }) === 5'b11000);
assign rom_instr_pt[22] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[2] , rom_addr_l2[4] ,
    rom_addr_l2[5] , rom_addr_l2[6] ,
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 8'b01101100);
assign rom_instr_pt[23] =
    (({ rom_addr_l2[1] , rom_addr_l2[4] ,
    rom_addr_l2[5] , rom_addr_l2[6] ,
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 6'b101100);
assign rom_instr_pt[24] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[2] , rom_addr_l2[6] ,
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 6'b010100);
assign rom_instr_pt[25] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] ,
    rom_addr_l2[3] , rom_addr_l2[5] ,
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 6'b000000);
assign rom_instr_pt[26] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[2] , rom_addr_l2[3] ,
    rom_addr_l2[5] , rom_addr_l2[7] ,
    rom_addr_l2[8] }) === 7'b0100000);
assign rom_instr_pt[27] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] ,
    rom_addr_l2[3] , rom_addr_l2[4] ,
    rom_addr_l2[5] , rom_addr_l2[7] ,
    rom_addr_l2[8] }) === 7'b0000100);
assign rom_instr_pt[28] =
    (({ rom_addr_l2[0] , rom_addr_l2[2] ,
    rom_addr_l2[3] , rom_addr_l2[4] ,
    rom_addr_l2[5] , rom_addr_l2[7] ,
    rom_addr_l2[8] }) === 7'b0001100);
assign rom_instr_pt[29] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[3] , rom_addr_l2[4] ,
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 6'b010100);
assign rom_instr_pt[30] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[2] , rom_addr_l2[3] ,
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 6'b010000);
assign rom_instr_pt[31] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[2] , rom_addr_l2[4] ,
    rom_addr_l2[5] , rom_addr_l2[6] ,
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 8'b01011010);
assign rom_instr_pt[32] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] ,
    rom_addr_l2[4] , rom_addr_l2[6] ,
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 6'b011010);
assign rom_instr_pt[33] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] ,
    rom_addr_l2[3] , rom_addr_l2[6] ,
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 6'b011010);
assign rom_instr_pt[34] =
    (({ rom_addr_l2[1] , rom_addr_l2[3] ,
    rom_addr_l2[6] , rom_addr_l2[7] ,
    rom_addr_l2[8] }) === 5'b10110);
assign rom_instr_pt[35] =
    (({ rom_addr_l2[3] , rom_addr_l2[6] ,
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 4'b0110);
assign rom_instr_pt[36] =
    (({ rom_addr_l2[1] , rom_addr_l2[3] ,
    rom_addr_l2[6] , rom_addr_l2[7] ,
    rom_addr_l2[8] }) === 5'b01110);
assign rom_instr_pt[37] =
    (({ rom_addr_l2[3] , rom_addr_l2[6] ,
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 4'b1110);
assign rom_instr_pt[38] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[3] , rom_addr_l2[4] ,
    rom_addr_l2[5] , rom_addr_l2[7] ,
    rom_addr_l2[8] }) === 7'b0110010);
assign rom_instr_pt[39] =
    (({ rom_addr_l2[1] , rom_addr_l2[4] ,
    rom_addr_l2[5] , rom_addr_l2[7] ,
    rom_addr_l2[8] }) === 5'b11010);
assign rom_instr_pt[40] =
    (({ rom_addr_l2[1] , rom_addr_l2[5] ,
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 4'b0010);
assign rom_instr_pt[41] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[2] , rom_addr_l2[3] ,
    rom_addr_l2[4] , rom_addr_l2[5] ,
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 8'b01010110);
assign rom_instr_pt[42] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[2] , rom_addr_l2[3] ,
    rom_addr_l2[5] , rom_addr_l2[7] ,
    rom_addr_l2[8] }) === 7'b0000110);
assign rom_instr_pt[43] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] ,
    rom_addr_l2[3] , rom_addr_l2[4] ,
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 6'b010010);
assign rom_instr_pt[44] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] ,
    rom_addr_l2[3] , rom_addr_l2[4] ,
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 6'b110010);
assign rom_instr_pt[45] =
    (({ rom_addr_l2[3] , rom_addr_l2[4] ,
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 4'b0010);
assign rom_instr_pt[46] =
    (({ rom_addr_l2[2] , rom_addr_l2[3] ,
    rom_addr_l2[4] , rom_addr_l2[7] ,
    rom_addr_l2[8] }) === 5'b11110);
assign rom_instr_pt[47] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[2] , rom_addr_l2[3] ,
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 6'b000010);
assign rom_instr_pt[48] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[2] , rom_addr_l2[3] ,
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 6'b010010);
assign rom_instr_pt[49] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] ,
    rom_addr_l2[3] , rom_addr_l2[7] ,
    rom_addr_l2[8] }) === 5'b00110);
assign rom_instr_pt[50] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[2] , rom_addr_l2[7] ,
    rom_addr_l2[8] }) === 5'b11010);
assign rom_instr_pt[51] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 4'b1010);
assign rom_instr_pt[52] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 4'b1110);
assign rom_instr_pt[53] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[2] , rom_addr_l2[3] ,
    rom_addr_l2[4] , rom_addr_l2[6] ,
    rom_addr_l2[8] }) === 7'b0111000);
assign rom_instr_pt[54] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[2] , rom_addr_l2[3] ,
    rom_addr_l2[6] , rom_addr_l2[8]
     }) === 6'b111000);
assign rom_instr_pt[55] =
    (({ rom_addr_l2[2] , rom_addr_l2[3] ,
    rom_addr_l2[4] , rom_addr_l2[6] ,
    rom_addr_l2[8] }) === 5'b10010);
assign rom_instr_pt[56] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[3] , rom_addr_l2[4] ,
    rom_addr_l2[6] , rom_addr_l2[8]
     }) === 6'b000010);
assign rom_instr_pt[57] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[3] , rom_addr_l2[4] ,
    rom_addr_l2[6] , rom_addr_l2[8]
     }) === 6'b100010);
assign rom_instr_pt[58] =
    (({ rom_addr_l2[1] , rom_addr_l2[3] ,
    rom_addr_l2[4] , rom_addr_l2[6] ,
    rom_addr_l2[8] }) === 5'b00010);
assign rom_instr_pt[59] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[2] , rom_addr_l2[4] ,
    rom_addr_l2[6] , rom_addr_l2[8]
     }) === 6'b100010);
assign rom_instr_pt[60] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[2] , rom_addr_l2[4] ,
    rom_addr_l2[6] , rom_addr_l2[8]
     }) === 6'b000110);
assign rom_instr_pt[61] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[2] , rom_addr_l2[3] ,
    rom_addr_l2[6] , rom_addr_l2[8]
     }) === 6'b111010);
assign rom_instr_pt[62] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[3] , rom_addr_l2[6] ,
    rom_addr_l2[8] }) === 5'b10110);
assign rom_instr_pt[63] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[2] , rom_addr_l2[6] ,
    rom_addr_l2[8] }) === 5'b00010);
assign rom_instr_pt[64] =
    (({ rom_addr_l2[1] , rom_addr_l2[5] ,
    rom_addr_l2[8] }) === 3'b000);
assign rom_instr_pt[65] =
    (({ rom_addr_l2[1] , rom_addr_l2[3] ,
    rom_addr_l2[4] , rom_addr_l2[8]
     }) === 4'b0000);
assign rom_instr_pt[66] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[3] , rom_addr_l2[4] ,
    rom_addr_l2[8] }) === 5'b01010);
assign rom_instr_pt[67] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[2] , rom_addr_l2[4] ,
    rom_addr_l2[8] }) === 5'b00110);
assign rom_instr_pt[68] =
    (({ rom_addr_l2[3] , rom_addr_l2[8]
     }) === 2'b00);
assign rom_instr_pt[69] =
    (({ rom_addr_l2[2] , rom_addr_l2[8]
     }) === 2'b00);
assign rom_instr_pt[70] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] ,
    rom_addr_l2[5] , rom_addr_l2[6] ,
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 6'b101001);
assign rom_instr_pt[71] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] ,
    rom_addr_l2[3] , rom_addr_l2[4] ,
    rom_addr_l2[6] , rom_addr_l2[7] ,
    rom_addr_l2[8] }) === 7'b0100001);
assign rom_instr_pt[72] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] ,
    rom_addr_l2[3] , rom_addr_l2[4] ,
    rom_addr_l2[6] , rom_addr_l2[7] ,
    rom_addr_l2[8] }) === 7'b1100001);
assign rom_instr_pt[73] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] ,
    rom_addr_l2[3] , rom_addr_l2[6] ,
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 6'b001001);
assign rom_instr_pt[74] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[6] , rom_addr_l2[7] ,
    rom_addr_l2[8] }) === 5'b11001);
assign rom_instr_pt[75] =
    (({ rom_addr_l2[2] , rom_addr_l2[4] ,
    rom_addr_l2[6] , rom_addr_l2[7] ,
    rom_addr_l2[8] }) === 5'b11101);
assign rom_instr_pt[76] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] ,
    rom_addr_l2[3] , rom_addr_l2[6] ,
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 6'b011101);
assign rom_instr_pt[77] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] ,
    rom_addr_l2[4] , rom_addr_l2[5] ,
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 6'b101001);
assign rom_instr_pt[78] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] ,
    rom_addr_l2[3] , rom_addr_l2[5] ,
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 6'b000001);
assign rom_instr_pt[79] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] ,
    rom_addr_l2[3] , rom_addr_l2[4] ,
    rom_addr_l2[5] , rom_addr_l2[7] ,
    rom_addr_l2[8] }) === 7'b0000101);
assign rom_instr_pt[80] =
    (({ rom_addr_l2[0] , rom_addr_l2[2] ,
    rom_addr_l2[3] , rom_addr_l2[4] ,
    rom_addr_l2[5] , rom_addr_l2[7] ,
    rom_addr_l2[8] }) === 7'b0001101);
assign rom_instr_pt[81] =
    (({ rom_addr_l2[2] , rom_addr_l2[3] ,
    rom_addr_l2[4] , rom_addr_l2[5] ,
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 6'b111101);
assign rom_instr_pt[82] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] ,
    rom_addr_l2[4] , rom_addr_l2[5] ,
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 6'b011101);
assign rom_instr_pt[83] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[3] , rom_addr_l2[4] ,
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 6'b010001);
assign rom_instr_pt[84] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[2] , rom_addr_l2[3] ,
    rom_addr_l2[4] , rom_addr_l2[7] ,
    rom_addr_l2[8] }) === 7'b0101001);
assign rom_instr_pt[85] =
    (({ rom_addr_l2[3] , rom_addr_l2[4] ,
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 4'b0101);
assign rom_instr_pt[86] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[4] , rom_addr_l2[7] ,
    rom_addr_l2[8] }) === 5'b10101);
assign rom_instr_pt[87] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[2] , rom_addr_l2[3] ,
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 6'b010001);
assign rom_instr_pt[88] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] ,
    rom_addr_l2[3] , rom_addr_l2[7] ,
    rom_addr_l2[8] }) === 5'b01101);
assign rom_instr_pt[89] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[2] , rom_addr_l2[7] ,
    rom_addr_l2[8] }) === 5'b11001);
assign rom_instr_pt[90] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[3] , rom_addr_l2[4] ,
    rom_addr_l2[6] , rom_addr_l2[7] ,
    rom_addr_l2[8] }) === 7'b0101011);
assign rom_instr_pt[91] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] ,
    rom_addr_l2[4] , rom_addr_l2[6] ,
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 6'b011011);
assign rom_instr_pt[92] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] ,
    rom_addr_l2[3] , rom_addr_l2[6] ,
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 6'b011011);
assign rom_instr_pt[93] =
    (({ rom_addr_l2[1] , rom_addr_l2[3] ,
    rom_addr_l2[6] , rom_addr_l2[7] ,
    rom_addr_l2[8] }) === 5'b11111);
assign rom_instr_pt[94] =
    (({ rom_addr_l2[3] , rom_addr_l2[6] ,
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 4'b1111);
assign rom_instr_pt[95] =
    (({ rom_addr_l2[1] , rom_addr_l2[4] ,
    rom_addr_l2[5] , rom_addr_l2[7] ,
    rom_addr_l2[8] }) === 5'b11011);
assign rom_instr_pt[96] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] ,
    rom_addr_l2[3] , rom_addr_l2[5] ,
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 6'b000011);
assign rom_instr_pt[97] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] ,
    rom_addr_l2[3] , rom_addr_l2[5] ,
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 6'b100011);
assign rom_instr_pt[98] =
    (({ rom_addr_l2[2] , rom_addr_l2[3] ,
    rom_addr_l2[5] , rom_addr_l2[7] ,
    rom_addr_l2[8] }) === 5'b00011);
assign rom_instr_pt[99] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[2] , rom_addr_l2[5] ,
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 6'b111011);
assign rom_instr_pt[100] =
    (({ rom_addr_l2[0] , rom_addr_l2[2] ,
    rom_addr_l2[3] , rom_addr_l2[4] ,
    rom_addr_l2[5] , rom_addr_l2[7] ,
    rom_addr_l2[8] }) === 7'b0001111);
assign rom_instr_pt[101] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[2] , rom_addr_l2[3] ,
    rom_addr_l2[5] , rom_addr_l2[7] ,
    rom_addr_l2[8] }) === 7'b0000111);
assign rom_instr_pt[102] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[2] , rom_addr_l2[3] ,
    rom_addr_l2[5] , rom_addr_l2[7] ,
    rom_addr_l2[8] }) === 7'b0100111);
assign rom_instr_pt[103] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[2] , rom_addr_l2[5] ,
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 6'b111111);
assign rom_instr_pt[104] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] ,
    rom_addr_l2[3] , rom_addr_l2[4] ,
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 6'b010011);
assign rom_instr_pt[105] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[2] , rom_addr_l2[3] ,
    rom_addr_l2[4] , rom_addr_l2[7] ,
    rom_addr_l2[8] }) === 7'b0101011);
assign rom_instr_pt[106] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[2] , rom_addr_l2[4] ,
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 6'b011011);
assign rom_instr_pt[107] =
    (({ rom_addr_l2[2] , rom_addr_l2[3] ,
    rom_addr_l2[4] , rom_addr_l2[7] ,
    rom_addr_l2[8] }) === 5'b11111);
assign rom_instr_pt[108] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[2] , rom_addr_l2[4] ,
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 6'b010111);
assign rom_instr_pt[109] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[2] , rom_addr_l2[3] ,
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 6'b000011);
assign rom_instr_pt[110] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] ,
    rom_addr_l2[3] , rom_addr_l2[7] ,
    rom_addr_l2[8] }) === 5'b10011);
assign rom_instr_pt[111] =
    (({ rom_addr_l2[2] , rom_addr_l2[3] ,
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 4'b0011);
assign rom_instr_pt[112] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] ,
    rom_addr_l2[3] , rom_addr_l2[7] ,
    rom_addr_l2[8] }) === 5'b00111);
assign rom_instr_pt[113] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[2] , rom_addr_l2[7] ,
    rom_addr_l2[8] }) === 5'b10011);
assign rom_instr_pt[114] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[2] , rom_addr_l2[7] ,
    rom_addr_l2[8] }) === 5'b11011);
assign rom_instr_pt[115] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] ,
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 4'b0111);
assign rom_instr_pt[116] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[2] , rom_addr_l2[7] ,
    rom_addr_l2[8] }) === 5'b11111);
assign rom_instr_pt[117] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[7] , rom_addr_l2[8]
     }) === 4'b1011);
assign rom_instr_pt[118] =
    (({ rom_addr_l2[2] , rom_addr_l2[4] ,
    rom_addr_l2[6] , rom_addr_l2[8]
     }) === 4'b1001);
assign rom_instr_pt[119] =
    (({ rom_addr_l2[0] , rom_addr_l2[5] ,
    rom_addr_l2[6] , rom_addr_l2[8]
     }) === 4'b1011);
assign rom_instr_pt[120] =
    (({ rom_addr_l2[5] , rom_addr_l2[6] ,
    rom_addr_l2[8] }) === 3'b011);
assign rom_instr_pt[121] =
    (({ rom_addr_l2[1] , rom_addr_l2[3] ,
    rom_addr_l2[4] , rom_addr_l2[5] ,
    rom_addr_l2[6] , rom_addr_l2[8]
     }) === 6'b000111);
assign rom_instr_pt[122] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[5] , rom_addr_l2[6] ,
    rom_addr_l2[8] }) === 5'b11111);
assign rom_instr_pt[123] =
    (({ rom_addr_l2[3] , rom_addr_l2[4] ,
    rom_addr_l2[6] , rom_addr_l2[8]
     }) === 4'b0011);
assign rom_instr_pt[124] =
    (({ rom_addr_l2[1] , rom_addr_l2[3] ,
    rom_addr_l2[4] , rom_addr_l2[6] ,
    rom_addr_l2[8] }) === 5'b11111);
assign rom_instr_pt[125] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] ,
    rom_addr_l2[4] , rom_addr_l2[6] ,
    rom_addr_l2[8] }) === 5'b01111);
assign rom_instr_pt[126] =
    (({ rom_addr_l2[1] , rom_addr_l2[3] ,
    rom_addr_l2[6] , rom_addr_l2[8]
     }) === 4'b0011);
assign rom_instr_pt[127] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] ,
    rom_addr_l2[3] , rom_addr_l2[6] ,
    rom_addr_l2[8] }) === 5'b11111);
assign rom_instr_pt[128] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] ,
    rom_addr_l2[6] , rom_addr_l2[8]
     }) === 4'b0011);
assign rom_instr_pt[129] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[6] , rom_addr_l2[8]
     }) === 4'b1111);
assign rom_instr_pt[130] =
    (({ rom_addr_l2[2] , rom_addr_l2[4] ,
    rom_addr_l2[5] , rom_addr_l2[8]
     }) === 4'b1101);
assign rom_instr_pt[131] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] ,
    rom_addr_l2[3] , rom_addr_l2[5] ,
    rom_addr_l2[8] }) === 5'b11101);
assign rom_instr_pt[132] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] ,
    rom_addr_l2[3] , rom_addr_l2[4] ,
    rom_addr_l2[5] , rom_addr_l2[8]
     }) === 6'b000011);
assign rom_instr_pt[133] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] ,
    rom_addr_l2[3] , rom_addr_l2[4] ,
    rom_addr_l2[8] }) === 5'b01111);
assign rom_instr_pt[134] =
    (({ rom_addr_l2[3] , rom_addr_l2[4] ,
    rom_addr_l2[8] }) === 3'b111);
assign rom_instr_pt[135] =
    (({ rom_addr_l2[1] , rom_addr_l2[3] ,
    rom_addr_l2[8] }) === 3'b011);
assign rom_instr_pt[136] =
    (({ rom_addr_l2[1] , rom_addr_l2[3] ,
    rom_addr_l2[4] , rom_addr_l2[5] ,
    rom_addr_l2[6] , rom_addr_l2[7]
     }) === 6'b000000);
assign rom_instr_pt[137] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] ,
    rom_addr_l2[5] , rom_addr_l2[6] ,
    rom_addr_l2[7] }) === 5'b00000);
assign rom_instr_pt[138] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[2] , rom_addr_l2[3] ,
    rom_addr_l2[4] , rom_addr_l2[6] ,
    rom_addr_l2[7] }) === 7'b0101000);
assign rom_instr_pt[139] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[2] , rom_addr_l2[3] ,
    rom_addr_l2[4] , rom_addr_l2[6] ,
    rom_addr_l2[7] }) === 7'b0111000);
assign rom_instr_pt[140] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] ,
    rom_addr_l2[3] , rom_addr_l2[4] ,
    rom_addr_l2[6] , rom_addr_l2[7]
     }) === 6'b111000);
assign rom_instr_pt[141] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] ,
    rom_addr_l2[3] , rom_addr_l2[6] ,
    rom_addr_l2[7] }) === 5'b01100);
assign rom_instr_pt[142] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[4] , rom_addr_l2[6] ,
    rom_addr_l2[7] }) === 5'b00110);
assign rom_instr_pt[143] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[2] , rom_addr_l2[3] ,
    rom_addr_l2[6] , rom_addr_l2[7]
     }) === 6'b001110);
assign rom_instr_pt[144] =
    (({ rom_addr_l2[0] , rom_addr_l2[2] ,
    rom_addr_l2[3] , rom_addr_l2[6] ,
    rom_addr_l2[7] }) === 5'b01110);
assign rom_instr_pt[145] =
    (({ rom_addr_l2[6] , rom_addr_l2[7]
     }) === 2'b10);
assign rom_instr_pt[146] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] ,
    rom_addr_l2[3] , rom_addr_l2[4] ,
    rom_addr_l2[5] , rom_addr_l2[7]
     }) === 6'b000010);
assign rom_instr_pt[147] =
    (({ rom_addr_l2[3] , rom_addr_l2[7]
     }) === 2'b00);
assign rom_instr_pt[148] =
    (({ rom_addr_l2[3] , rom_addr_l2[4] ,
    rom_addr_l2[6] , rom_addr_l2[7]
     }) === 4'b1111);
assign rom_instr_pt[149] =
    (({ rom_addr_l2[1] , rom_addr_l2[6] ,
    rom_addr_l2[7] }) === 3'b111);
assign rom_instr_pt[150] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] ,
    rom_addr_l2[4] , rom_addr_l2[5] ,
    rom_addr_l2[7] }) === 5'b11011);
assign rom_instr_pt[151] =
    (({ rom_addr_l2[2] , rom_addr_l2[4] ,
    rom_addr_l2[7] }) === 3'b011);
assign rom_instr_pt[152] =
    (({ rom_addr_l2[2] , rom_addr_l2[3] ,
    rom_addr_l2[7] }) === 3'b011);
assign rom_instr_pt[153] =
    (({ rom_addr_l2[2] , rom_addr_l2[3] ,
    rom_addr_l2[4] , rom_addr_l2[5] ,
    rom_addr_l2[6] }) === 5'b10100);
assign rom_instr_pt[154] =
    (({ rom_addr_l2[0] , rom_addr_l2[2] ,
    rom_addr_l2[3] , rom_addr_l2[5] ,
    rom_addr_l2[6] }) === 5'b11100);
assign rom_instr_pt[155] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[3] , rom_addr_l2[4] ,
    rom_addr_l2[5] , rom_addr_l2[6]
     }) === 6'b010110);
assign rom_instr_pt[156] =
    (({ rom_addr_l2[0] , rom_addr_l2[2] ,
    rom_addr_l2[3] , rom_addr_l2[4] ,
    rom_addr_l2[6] }) === 5'b10000);
assign rom_instr_pt[157] =
    (({ rom_addr_l2[0] , rom_addr_l2[3] ,
    rom_addr_l2[4] , rom_addr_l2[6]
     }) === 4'b0010);
assign rom_instr_pt[158] =
    (({ rom_addr_l2[0] , rom_addr_l2[2] ,
    rom_addr_l2[4] , rom_addr_l2[6]
     }) === 4'b1010);
assign rom_instr_pt[159] =
    (({ rom_addr_l2[0] , rom_addr_l2[2] ,
    rom_addr_l2[4] , rom_addr_l2[6]
     }) === 4'b1110);
assign rom_instr_pt[160] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[2] , rom_addr_l2[3] ,
    rom_addr_l2[6] }) === 5'b11100);
assign rom_instr_pt[161] =
    (({ rom_addr_l2[2] , rom_addr_l2[3] ,
    rom_addr_l2[6] }) === 3'b010);
assign rom_instr_pt[162] =
    (({ rom_addr_l2[0] , rom_addr_l2[2] ,
    rom_addr_l2[3] , rom_addr_l2[6]
     }) === 4'b1110);
assign rom_instr_pt[163] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[2] , rom_addr_l2[4] ,
    rom_addr_l2[5] , rom_addr_l2[6]
     }) === 6'b010001);
assign rom_instr_pt[164] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[4] , rom_addr_l2[5] ,
    rom_addr_l2[6] }) === 5'b00101);
assign rom_instr_pt[165] =
    (({ rom_addr_l2[1] , rom_addr_l2[4] ,
    rom_addr_l2[5] , rom_addr_l2[6]
     }) === 4'b1101);
assign rom_instr_pt[166] =
    (({ rom_addr_l2[0] , rom_addr_l2[4] ,
    rom_addr_l2[5] , rom_addr_l2[6]
     }) === 4'b1101);
assign rom_instr_pt[167] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[2] , rom_addr_l2[5] ,
    rom_addr_l2[6] }) === 5'b11001);
assign rom_instr_pt[168] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[2] , rom_addr_l2[5] ,
    rom_addr_l2[6] }) === 5'b01101);
assign rom_instr_pt[169] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[2] , rom_addr_l2[4] ,
    rom_addr_l2[5] , rom_addr_l2[6]
     }) === 6'b010011);
assign rom_instr_pt[170] =
    (({ rom_addr_l2[0] , rom_addr_l2[3] ,
    rom_addr_l2[4] , rom_addr_l2[5] ,
    rom_addr_l2[6] }) === 5'b11111);
assign rom_instr_pt[171] =
    (({ rom_addr_l2[0] , rom_addr_l2[2] ,
    rom_addr_l2[4] , rom_addr_l2[5] ,
    rom_addr_l2[6] }) === 5'b11111);
assign rom_instr_pt[172] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[3] , rom_addr_l2[5] ,
    rom_addr_l2[6] }) === 5'b10111);
assign rom_instr_pt[173] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[2] , rom_addr_l2[5] ,
    rom_addr_l2[6] }) === 5'b11011);
assign rom_instr_pt[174] =
    (({ rom_addr_l2[2] , rom_addr_l2[3] ,
    rom_addr_l2[4] , rom_addr_l2[6]
     }) === 4'b0001);
assign rom_instr_pt[175] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[2] , rom_addr_l2[4] ,
    rom_addr_l2[6] }) === 5'b01001);
assign rom_instr_pt[176] =
    (({ rom_addr_l2[4] , rom_addr_l2[6]
     }) === 2'b01);
assign rom_instr_pt[177] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[2] , rom_addr_l2[4] ,
    rom_addr_l2[6] }) === 5'b10011);
assign rom_instr_pt[178] =
    (({ rom_addr_l2[0] , rom_addr_l2[2] ,
    rom_addr_l2[4] , rom_addr_l2[6]
     }) === 4'b1011);
assign rom_instr_pt[179] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[4] , rom_addr_l2[6]
     }) === 4'b1011);
assign rom_instr_pt[180] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[2] , rom_addr_l2[3] ,
    rom_addr_l2[6] }) === 5'b11111);
assign rom_instr_pt[181] =
    (({ rom_addr_l2[0] , rom_addr_l2[2] ,
    rom_addr_l2[3] , rom_addr_l2[6]
     }) === 4'b1111);
assign rom_instr_pt[182] =
    (({ rom_addr_l2[0] , rom_addr_l2[3] ,
    rom_addr_l2[6] }) === 3'b111);
assign rom_instr_pt[183] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[2] , rom_addr_l2[6]
     }) === 4'b0001);
assign rom_instr_pt[184] =
    (({ rom_addr_l2[2] , rom_addr_l2[6]
     }) === 2'b01);
assign rom_instr_pt[185] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[2] , rom_addr_l2[6]
     }) === 4'b0111);
assign rom_instr_pt[186] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[6] }) === 3'b011);
assign rom_instr_pt[187] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[2] , rom_addr_l2[3] ,
    rom_addr_l2[4] , rom_addr_l2[5]
     }) === 6'b001100);
assign rom_instr_pt[188] =
    (({ rom_addr_l2[1] , rom_addr_l2[4] ,
    rom_addr_l2[5] }) === 3'b000);
assign rom_instr_pt[189] =
    (({ rom_addr_l2[1] , rom_addr_l2[3] ,
    rom_addr_l2[4] , rom_addr_l2[5]
     }) === 4'b1110);
assign rom_instr_pt[190] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] ,
    rom_addr_l2[3] , rom_addr_l2[4] ,
    rom_addr_l2[5] }) === 5'b01001);
assign rom_instr_pt[191] =
    (({ rom_addr_l2[2] , rom_addr_l2[3] ,
    rom_addr_l2[4] , rom_addr_l2[5]
     }) === 4'b1111);
assign rom_instr_pt[192] =
    (({ rom_addr_l2[0] , rom_addr_l2[1] ,
    rom_addr_l2[2] , rom_addr_l2[4] ,
    rom_addr_l2[5] }) === 5'b01011);
assign rom_instr_pt[193] =
    (({ rom_addr_l2[3] , rom_addr_l2[5]
     }) === 2'b11);
assign rom_instr_pt[194] =
    (({ rom_addr_l2[0] , rom_addr_l2[2] ,
    rom_addr_l2[3] , rom_addr_l2[4]
     }) === 4'b1000);
assign rom_instr_pt[195] =
    (({ rom_addr_l2[2] , rom_addr_l2[3] ,
    rom_addr_l2[4] }) === 3'b111);
assign rom_instr_pt[196] =
    (({ rom_addr_l2[3] , rom_addr_l2[4]
     }) === 2'b11);
assign rom_instr_pt[197] =
    (({ rom_addr_l2[1] , rom_addr_l2[4]
     }) === 2'b11);
assign rom_instr_pt[198] =
    (({ rom_addr_l2[1] , rom_addr_l2[2] ,
    rom_addr_l2[3] }) === 3'b001);
assign rom_instr_pt[199] =
    (({ rom_addr_l2[2] }) === 1'b0);
assign rom_instr_pt[200] =
    (({ rom_addr_l2[0] }) === 1'b1);
assign template[0] =
    (rom_instr_pt[1] | rom_instr_pt[4]
     | rom_instr_pt[25] | rom_instr_pt[29]
     | rom_instr_pt[38] | rom_instr_pt[80]
     | rom_instr_pt[99] | rom_instr_pt[155]
     | rom_instr_pt[166] | rom_instr_pt[167]
     | rom_instr_pt[168] | rom_instr_pt[171]
     | rom_instr_pt[181]);
assign template[1] =
    (rom_instr_pt[3] | rom_instr_pt[6]
     | rom_instr_pt[9] | rom_instr_pt[10]
     | rom_instr_pt[14] | rom_instr_pt[16]
     | rom_instr_pt[17] | rom_instr_pt[23]
     | rom_instr_pt[27] | rom_instr_pt[28]
     | rom_instr_pt[32] | rom_instr_pt[33]
     | rom_instr_pt[35] | rom_instr_pt[36]
     | rom_instr_pt[39] | rom_instr_pt[40]
     | rom_instr_pt[41] | rom_instr_pt[42]
     | rom_instr_pt[43] | rom_instr_pt[44]
     | rom_instr_pt[46] | rom_instr_pt[48]
     | rom_instr_pt[49] | rom_instr_pt[50]
     | rom_instr_pt[51] | rom_instr_pt[53]
     | rom_instr_pt[54] | rom_instr_pt[57]
     | rom_instr_pt[59] | rom_instr_pt[61]
     | rom_instr_pt[71] | rom_instr_pt[72]
     | rom_instr_pt[73] | rom_instr_pt[76]
     | rom_instr_pt[78] | rom_instr_pt[82]
     | rom_instr_pt[84] | rom_instr_pt[86]
     | rom_instr_pt[87] | rom_instr_pt[89]
     | rom_instr_pt[91] | rom_instr_pt[92]
     | rom_instr_pt[94] | rom_instr_pt[103]
     | rom_instr_pt[104] | rom_instr_pt[105]
     | rom_instr_pt[109] | rom_instr_pt[112]
     | rom_instr_pt[113] | rom_instr_pt[122]
     | rom_instr_pt[125] | rom_instr_pt[127]
     | rom_instr_pt[132] | rom_instr_pt[134]
     | rom_instr_pt[139] | rom_instr_pt[165]
     | rom_instr_pt[172] | rom_instr_pt[173]
     | rom_instr_pt[177] | rom_instr_pt[180]
     | rom_instr_pt[183] | rom_instr_pt[192]
     | rom_instr_pt[194]);
assign template[2] =
    (rom_instr_pt[6] | rom_instr_pt[8]
     | rom_instr_pt[10] | rom_instr_pt[17]
     | rom_instr_pt[19] | rom_instr_pt[21]
     | rom_instr_pt[22] | rom_instr_pt[24]
     | rom_instr_pt[27] | rom_instr_pt[28]
     | rom_instr_pt[33] | rom_instr_pt[36]
     | rom_instr_pt[40] | rom_instr_pt[41]
     | rom_instr_pt[43] | rom_instr_pt[44]
     | rom_instr_pt[49] | rom_instr_pt[51]
     | rom_instr_pt[56] | rom_instr_pt[57]
     | rom_instr_pt[59] | rom_instr_pt[61]
     | rom_instr_pt[71] | rom_instr_pt[72]
     | rom_instr_pt[103] | rom_instr_pt[104]
     | rom_instr_pt[106] | rom_instr_pt[109]
     | rom_instr_pt[110] | rom_instr_pt[114]
     | rom_instr_pt[123] | rom_instr_pt[125]
     | rom_instr_pt[132] | rom_instr_pt[139]
     | rom_instr_pt[141] | rom_instr_pt[142]
     | rom_instr_pt[143] | rom_instr_pt[149]
     | rom_instr_pt[153] | rom_instr_pt[171]
     | rom_instr_pt[172] | rom_instr_pt[173]
     | rom_instr_pt[177] | rom_instr_pt[183]
     | rom_instr_pt[192] | rom_instr_pt[194]
     | rom_instr_pt[195]);
assign template[3] =
    (rom_instr_pt[3] | rom_instr_pt[6]
     | rom_instr_pt[8] | rom_instr_pt[10]
     | rom_instr_pt[14] | rom_instr_pt[17]
     | rom_instr_pt[19] | rom_instr_pt[20]
     | rom_instr_pt[21] | rom_instr_pt[22]
     | rom_instr_pt[24] | rom_instr_pt[27]
     | rom_instr_pt[28] | rom_instr_pt[29]
     | rom_instr_pt[32] | rom_instr_pt[33]
     | rom_instr_pt[35] | rom_instr_pt[36]
     | rom_instr_pt[38] | rom_instr_pt[39]
     | rom_instr_pt[40] | rom_instr_pt[41]
     | rom_instr_pt[42] | rom_instr_pt[43]
     | rom_instr_pt[44] | rom_instr_pt[46]
     | rom_instr_pt[48] | rom_instr_pt[49]
     | rom_instr_pt[50] | rom_instr_pt[51]
     | rom_instr_pt[53] | rom_instr_pt[56]
     | rom_instr_pt[59] | rom_instr_pt[61]
     | rom_instr_pt[71] | rom_instr_pt[72]
     | rom_instr_pt[73] | rom_instr_pt[77]
     | rom_instr_pt[78] | rom_instr_pt[79]
     | rom_instr_pt[81] | rom_instr_pt[82]
     | rom_instr_pt[84] | rom_instr_pt[86]
     | rom_instr_pt[87] | rom_instr_pt[89]
     | rom_instr_pt[91] | rom_instr_pt[92]
     | rom_instr_pt[94] | rom_instr_pt[95]
     | rom_instr_pt[99] | rom_instr_pt[100]
     | rom_instr_pt[103] | rom_instr_pt[104]
     | rom_instr_pt[105] | rom_instr_pt[106]
     | rom_instr_pt[107] | rom_instr_pt[110]
     | rom_instr_pt[112] | rom_instr_pt[113]
     | rom_instr_pt[114] | rom_instr_pt[123]
     | rom_instr_pt[125] | rom_instr_pt[127]
     | rom_instr_pt[128] | rom_instr_pt[139]
     | rom_instr_pt[141] | rom_instr_pt[142]
     | rom_instr_pt[143] | rom_instr_pt[149]
     | rom_instr_pt[153] | rom_instr_pt[155]
     | rom_instr_pt[167] | rom_instr_pt[168]
     | rom_instr_pt[173] | rom_instr_pt[177]
     | rom_instr_pt[192]);
assign template[4] =
    (rom_instr_pt[1] | rom_instr_pt[4]
     | rom_instr_pt[6] | rom_instr_pt[8]
     | rom_instr_pt[10] | rom_instr_pt[17]
     | rom_instr_pt[19] | rom_instr_pt[20]
     | rom_instr_pt[21] | rom_instr_pt[23]
     | rom_instr_pt[24] | rom_instr_pt[25]
     | rom_instr_pt[27] | rom_instr_pt[28]
     | rom_instr_pt[29] | rom_instr_pt[33]
     | rom_instr_pt[36] | rom_instr_pt[38]
     | rom_instr_pt[40] | rom_instr_pt[41]
     | rom_instr_pt[43] | rom_instr_pt[44]
     | rom_instr_pt[46] | rom_instr_pt[49]
     | rom_instr_pt[51] | rom_instr_pt[56]
     | rom_instr_pt[57] | rom_instr_pt[59]
     | rom_instr_pt[61] | rom_instr_pt[71]
     | rom_instr_pt[72] | rom_instr_pt[80]
     | rom_instr_pt[81] | rom_instr_pt[99]
     | rom_instr_pt[103] | rom_instr_pt[104]
     | rom_instr_pt[106] | rom_instr_pt[107]
     | rom_instr_pt[109] | rom_instr_pt[110]
     | rom_instr_pt[114] | rom_instr_pt[123]
     | rom_instr_pt[125] | rom_instr_pt[132]
     | rom_instr_pt[139] | rom_instr_pt[141]
     | rom_instr_pt[142] | rom_instr_pt[143]
     | rom_instr_pt[149] | rom_instr_pt[153]
     | rom_instr_pt[155] | rom_instr_pt[166]
     | rom_instr_pt[167] | rom_instr_pt[168]
     | rom_instr_pt[172] | rom_instr_pt[173]
     | rom_instr_pt[177] | rom_instr_pt[183]
     | rom_instr_pt[192]);
assign template[5] =
    (rom_instr_pt[3] | rom_instr_pt[6]
     | rom_instr_pt[9] | rom_instr_pt[10]
     | rom_instr_pt[14] | rom_instr_pt[16]
     | rom_instr_pt[17] | rom_instr_pt[22]
     | rom_instr_pt[27] | rom_instr_pt[28]
     | rom_instr_pt[33] | rom_instr_pt[35]
     | rom_instr_pt[36] | rom_instr_pt[39]
     | rom_instr_pt[40] | rom_instr_pt[41]
     | rom_instr_pt[42] | rom_instr_pt[43]
     | rom_instr_pt[46] | rom_instr_pt[48]
     | rom_instr_pt[49] | rom_instr_pt[51]
     | rom_instr_pt[53] | rom_instr_pt[59]
     | rom_instr_pt[60] | rom_instr_pt[73]
     | rom_instr_pt[76] | rom_instr_pt[77]
     | rom_instr_pt[79] | rom_instr_pt[81]
     | rom_instr_pt[82] | rom_instr_pt[86]
     | rom_instr_pt[89] | rom_instr_pt[94]
     | rom_instr_pt[95] | rom_instr_pt[100]
     | rom_instr_pt[103] | rom_instr_pt[105]
     | rom_instr_pt[107] | rom_instr_pt[122]
     | rom_instr_pt[125] | rom_instr_pt[127]
     | rom_instr_pt[128] | rom_instr_pt[139]
     | rom_instr_pt[165] | rom_instr_pt[169]
     | rom_instr_pt[173] | rom_instr_pt[177]
     | rom_instr_pt[192] | rom_instr_pt[194]
    );
assign template[6] =
    1'b0;
assign template[7] =
    1'b0;
assign template[8] =
    1'b0;
assign template[9] =
    (rom_instr_pt[1] | rom_instr_pt[4]
     | rom_instr_pt[6] | rom_instr_pt[10]
     | rom_instr_pt[16] | rom_instr_pt[17]
     | rom_instr_pt[23] | rom_instr_pt[29]
     | rom_instr_pt[35] | rom_instr_pt[36]
     | rom_instr_pt[38] | rom_instr_pt[40]
     | rom_instr_pt[41] | rom_instr_pt[42]
     | rom_instr_pt[43] | rom_instr_pt[48]
     | rom_instr_pt[49] | rom_instr_pt[51]
     | rom_instr_pt[53] | rom_instr_pt[56]
     | rom_instr_pt[61] | rom_instr_pt[71]
     | rom_instr_pt[73] | rom_instr_pt[80]
     | rom_instr_pt[82] | rom_instr_pt[86]
     | rom_instr_pt[94] | rom_instr_pt[99]
     | rom_instr_pt[100] | rom_instr_pt[103]
     | rom_instr_pt[105] | rom_instr_pt[112]
     | rom_instr_pt[113] | rom_instr_pt[125]
     | rom_instr_pt[127] | rom_instr_pt[132]
     | rom_instr_pt[139] | rom_instr_pt[155]
     | rom_instr_pt[167] | rom_instr_pt[168]
     | rom_instr_pt[173] | rom_instr_pt[183]
    );
assign template[10] =
    (rom_instr_pt[25] | rom_instr_pt[27]
     | rom_instr_pt[32] | rom_instr_pt[33]
     | rom_instr_pt[39] | rom_instr_pt[44]
     | rom_instr_pt[50] | rom_instr_pt[54]
     | rom_instr_pt[57] | rom_instr_pt[72]
     | rom_instr_pt[76] | rom_instr_pt[77]
     | rom_instr_pt[78] | rom_instr_pt[89]
     | rom_instr_pt[91] | rom_instr_pt[92]
     | rom_instr_pt[95] | rom_instr_pt[104]
     | rom_instr_pt[121] | rom_instr_pt[165]
    );
assign template[11] =
    (rom_instr_pt[9] | rom_instr_pt[46]
     | rom_instr_pt[81] | rom_instr_pt[107]
     | rom_instr_pt[192]);
assign template[12] =
    1'b0;
assign template[13] =
    (rom_instr_pt[9]);
assign template[14] =
    (rom_instr_pt[14] | rom_instr_pt[16]
     | rom_instr_pt[32] | rom_instr_pt[35]
     | rom_instr_pt[40] | rom_instr_pt[42]
     | rom_instr_pt[43] | rom_instr_pt[44]
     | rom_instr_pt[48] | rom_instr_pt[49]
     | rom_instr_pt[50] | rom_instr_pt[51]
     | rom_instr_pt[53] | rom_instr_pt[54]
     | rom_instr_pt[57] | rom_instr_pt[61]
     | rom_instr_pt[70] | rom_instr_pt[71]
     | rom_instr_pt[73] | rom_instr_pt[78]
     | rom_instr_pt[82] | rom_instr_pt[84]
     | rom_instr_pt[86] | rom_instr_pt[87]
     | rom_instr_pt[89] | rom_instr_pt[91]
     | rom_instr_pt[92] | rom_instr_pt[94]
     | rom_instr_pt[105] | rom_instr_pt[112]
     | rom_instr_pt[113] | rom_instr_pt[125]
     | rom_instr_pt[127]);
assign template[15] =
    (rom_instr_pt[3] | rom_instr_pt[31]
     | rom_instr_pt[56] | rom_instr_pt[72]
     | rom_instr_pt[81] | rom_instr_pt[104]
     | rom_instr_pt[128]);
assign template[16] =
    (rom_instr_pt[32] | rom_instr_pt[39]
     | rom_instr_pt[50] | rom_instr_pt[77]
     | rom_instr_pt[82] | rom_instr_pt[84]
     | rom_instr_pt[92] | rom_instr_pt[108]
     | rom_instr_pt[112] | rom_instr_pt[113]
     | rom_instr_pt[121]);
assign template[17] =
    (rom_instr_pt[24] | rom_instr_pt[35]
     | rom_instr_pt[39] | rom_instr_pt[42]
     | rom_instr_pt[44] | rom_instr_pt[46]
     | rom_instr_pt[48] | rom_instr_pt[53]
     | rom_instr_pt[54] | rom_instr_pt[61]
     | rom_instr_pt[71] | rom_instr_pt[72]
     | rom_instr_pt[73] | rom_instr_pt[77]
     | rom_instr_pt[78] | rom_instr_pt[82]
     | rom_instr_pt[86] | rom_instr_pt[91]
     | rom_instr_pt[94] | rom_instr_pt[104]
     | rom_instr_pt[105] | rom_instr_pt[121]
     | rom_instr_pt[127]);
assign template[18] =
    (rom_instr_pt[77] | rom_instr_pt[121]
     | rom_instr_pt[124]);
assign template[19] =
    (rom_instr_pt[59] | rom_instr_pt[79]
     | rom_instr_pt[107] | rom_instr_pt[121]
     | rom_instr_pt[148] | rom_instr_pt[177]
    );
assign template[20] =
    (rom_instr_pt[16] | rom_instr_pt[36]
     | rom_instr_pt[40] | rom_instr_pt[43]
     | rom_instr_pt[49] | rom_instr_pt[51]
     | rom_instr_pt[79] | rom_instr_pt[121]
     | rom_instr_pt[125] | rom_instr_pt[194]
    );
assign template[21] =
    (rom_instr_pt[42] | rom_instr_pt[59]
     | rom_instr_pt[60] | rom_instr_pt[71]
     | rom_instr_pt[78] | rom_instr_pt[87]
     | rom_instr_pt[91] | rom_instr_pt[95]
     | rom_instr_pt[100] | rom_instr_pt[112]
     | rom_instr_pt[113] | rom_instr_pt[121]
     | rom_instr_pt[177]);
assign template[22] =
    (rom_instr_pt[16] | rom_instr_pt[28]
     | rom_instr_pt[32] | rom_instr_pt[36]
     | rom_instr_pt[39] | rom_instr_pt[40]
     | rom_instr_pt[43] | rom_instr_pt[49]
     | rom_instr_pt[51] | rom_instr_pt[60]
     | rom_instr_pt[87] | rom_instr_pt[92]
     | rom_instr_pt[100] | rom_instr_pt[123]
     | rom_instr_pt[125] | rom_instr_pt[128]
     | rom_instr_pt[169]);
assign template[23] =
    (rom_instr_pt[8] | rom_instr_pt[16]
     | rom_instr_pt[22] | rom_instr_pt[36]
     | rom_instr_pt[40] | rom_instr_pt[41]
     | rom_instr_pt[43] | rom_instr_pt[46]
     | rom_instr_pt[49] | rom_instr_pt[51]
     | rom_instr_pt[60] | rom_instr_pt[71]
     | rom_instr_pt[77] | rom_instr_pt[81]
     | rom_instr_pt[100] | rom_instr_pt[103]
     | rom_instr_pt[107] | rom_instr_pt[121]
     | rom_instr_pt[125] | rom_instr_pt[139]
     | rom_instr_pt[165] | rom_instr_pt[173]
    );
assign template[24] =
    (rom_instr_pt[6] | rom_instr_pt[10]
     | rom_instr_pt[17] | rom_instr_pt[22]
     | rom_instr_pt[27] | rom_instr_pt[33]
     | rom_instr_pt[41] | rom_instr_pt[59]
     | rom_instr_pt[60] | rom_instr_pt[71]
     | rom_instr_pt[76] | rom_instr_pt[79]
     | rom_instr_pt[103] | rom_instr_pt[121]
     | rom_instr_pt[139] | rom_instr_pt[173]
     | rom_instr_pt[177]);
assign template[25] =
    (rom_instr_pt[16] | rom_instr_pt[36]
     | rom_instr_pt[40] | rom_instr_pt[43]
     | rom_instr_pt[49] | rom_instr_pt[51]
     | rom_instr_pt[59] | rom_instr_pt[71]
     | rom_instr_pt[121] | rom_instr_pt[125]
     | rom_instr_pt[177]);
assign template[26] =
    (rom_instr_pt[6] | rom_instr_pt[9]
     | rom_instr_pt[10] | rom_instr_pt[14]
     | rom_instr_pt[16] | rom_instr_pt[17]
     | rom_instr_pt[22] | rom_instr_pt[27]
     | rom_instr_pt[33] | rom_instr_pt[35]
     | rom_instr_pt[36] | rom_instr_pt[39]
     | rom_instr_pt[40] | rom_instr_pt[41]
     | rom_instr_pt[42] | rom_instr_pt[43]
     | rom_instr_pt[46] | rom_instr_pt[48]
     | rom_instr_pt[49] | rom_instr_pt[51]
     | rom_instr_pt[53] | rom_instr_pt[59]
     | rom_instr_pt[60] | rom_instr_pt[71]
     | rom_instr_pt[73] | rom_instr_pt[76]
     | rom_instr_pt[77] | rom_instr_pt[78]
     | rom_instr_pt[79] | rom_instr_pt[81]
     | rom_instr_pt[82] | rom_instr_pt[86]
     | rom_instr_pt[87] | rom_instr_pt[89]
     | rom_instr_pt[91] | rom_instr_pt[94]
     | rom_instr_pt[95] | rom_instr_pt[100]
     | rom_instr_pt[103] | rom_instr_pt[105]
     | rom_instr_pt[107] | rom_instr_pt[112]
     | rom_instr_pt[113] | rom_instr_pt[121]
     | rom_instr_pt[125] | rom_instr_pt[127]
     | rom_instr_pt[139] | rom_instr_pt[165]
     | rom_instr_pt[173] | rom_instr_pt[177]
     | rom_instr_pt[192] | rom_instr_pt[194]
    );
assign template[27] =
    (rom_instr_pt[14] | rom_instr_pt[16]
     | rom_instr_pt[28] | rom_instr_pt[32]
     | rom_instr_pt[36] | rom_instr_pt[39]
     | rom_instr_pt[40] | rom_instr_pt[43]
     | rom_instr_pt[48] | rom_instr_pt[49]
     | rom_instr_pt[51] | rom_instr_pt[53]
     | rom_instr_pt[59] | rom_instr_pt[60]
     | rom_instr_pt[73] | rom_instr_pt[77]
     | rom_instr_pt[82] | rom_instr_pt[86]
     | rom_instr_pt[87] | rom_instr_pt[89]
     | rom_instr_pt[92] | rom_instr_pt[95]
     | rom_instr_pt[100] | rom_instr_pt[105]
     | rom_instr_pt[123] | rom_instr_pt[125]
     | rom_instr_pt[127] | rom_instr_pt[128]
     | rom_instr_pt[169] | rom_instr_pt[177]
    );
assign template[28] =
    (rom_instr_pt[6] | rom_instr_pt[10]
     | rom_instr_pt[14] | rom_instr_pt[16]
     | rom_instr_pt[17] | rom_instr_pt[22]
     | rom_instr_pt[27] | rom_instr_pt[32]
     | rom_instr_pt[33] | rom_instr_pt[35]
     | rom_instr_pt[36] | rom_instr_pt[39]
     | rom_instr_pt[40] | rom_instr_pt[41]
     | rom_instr_pt[42] | rom_instr_pt[43]
     | rom_instr_pt[48] | rom_instr_pt[49]
     | rom_instr_pt[50] | rom_instr_pt[51]
     | rom_instr_pt[53] | rom_instr_pt[59]
     | rom_instr_pt[73] | rom_instr_pt[76]
     | rom_instr_pt[77] | rom_instr_pt[78]
     | rom_instr_pt[79] | rom_instr_pt[82]
     | rom_instr_pt[84] | rom_instr_pt[86]
     | rom_instr_pt[87] | rom_instr_pt[89]
     | rom_instr_pt[91] | rom_instr_pt[92]
     | rom_instr_pt[94] | rom_instr_pt[95]
     | rom_instr_pt[103] | rom_instr_pt[105]
     | rom_instr_pt[112] | rom_instr_pt[113]
     | rom_instr_pt[121] | rom_instr_pt[125]
     | rom_instr_pt[127] | rom_instr_pt[139]
     | rom_instr_pt[173] | rom_instr_pt[177]
    );
assign template[29] =
    (rom_instr_pt[3] | rom_instr_pt[6]
     | rom_instr_pt[10] | rom_instr_pt[14]
     | rom_instr_pt[17] | rom_instr_pt[22]
     | rom_instr_pt[27] | rom_instr_pt[28]
     | rom_instr_pt[32] | rom_instr_pt[33]
     | rom_instr_pt[35] | rom_instr_pt[39]
     | rom_instr_pt[41] | rom_instr_pt[42]
     | rom_instr_pt[48] | rom_instr_pt[50]
     | rom_instr_pt[53] | rom_instr_pt[59]
     | rom_instr_pt[71] | rom_instr_pt[73]
     | rom_instr_pt[76] | rom_instr_pt[77]
     | rom_instr_pt[78] | rom_instr_pt[79]
     | rom_instr_pt[82] | rom_instr_pt[84]
     | rom_instr_pt[86] | rom_instr_pt[87]
     | rom_instr_pt[89] | rom_instr_pt[91]
     | rom_instr_pt[92] | rom_instr_pt[94]
     | rom_instr_pt[95] | rom_instr_pt[100]
     | rom_instr_pt[103] | rom_instr_pt[105]
     | rom_instr_pt[112] | rom_instr_pt[113]
     | rom_instr_pt[122] | rom_instr_pt[127]
     | rom_instr_pt[128] | rom_instr_pt[139]
     | rom_instr_pt[142] | rom_instr_pt[153]
     | rom_instr_pt[169] | rom_instr_pt[173]
     | rom_instr_pt[192]);
assign template[30] =
    (rom_instr_pt[3] | rom_instr_pt[6]
     | rom_instr_pt[10] | rom_instr_pt[14]
     | rom_instr_pt[17] | rom_instr_pt[22]
     | rom_instr_pt[27] | rom_instr_pt[29]
     | rom_instr_pt[32] | rom_instr_pt[33]
     | rom_instr_pt[35] | rom_instr_pt[39]
     | rom_instr_pt[41] | rom_instr_pt[42]
     | rom_instr_pt[48] | rom_instr_pt[50]
     | rom_instr_pt[53] | rom_instr_pt[73]
     | rom_instr_pt[76] | rom_instr_pt[77]
     | rom_instr_pt[78] | rom_instr_pt[79]
     | rom_instr_pt[82] | rom_instr_pt[84]
     | rom_instr_pt[86] | rom_instr_pt[87]
     | rom_instr_pt[89] | rom_instr_pt[90]
     | rom_instr_pt[91] | rom_instr_pt[92]
     | rom_instr_pt[94] | rom_instr_pt[95]
     | rom_instr_pt[103] | rom_instr_pt[105]
     | rom_instr_pt[112] | rom_instr_pt[113]
     | rom_instr_pt[127] | rom_instr_pt[139]
     | rom_instr_pt[170] | rom_instr_pt[173]
     | rom_instr_pt[192]);
assign template[31] =
    (rom_instr_pt[20] | rom_instr_pt[30]
     | rom_instr_pt[66] | rom_instr_pt[80]
     | rom_instr_pt[88] | rom_instr_pt[106]
     | rom_instr_pt[114] | rom_instr_pt[121]
     | rom_instr_pt[143] | rom_instr_pt[149]
    );
assign ucode_end =
    (rom_instr_pt[98] | rom_instr_pt[107]
     | rom_instr_pt[120] | rom_instr_pt[128]
     | rom_instr_pt[129] | rom_instr_pt[131]
     | rom_instr_pt[156] | rom_instr_pt[159]
     | rom_instr_pt[162] | rom_instr_pt[164]
     | rom_instr_pt[175] | rom_instr_pt[178]
    );
assign ucode_end_early =
    (rom_instr_pt[111] | rom_instr_pt[184]
     | rom_instr_pt[186]);
assign loop_begin =
    1'b0;
assign loop_end =
    (rom_instr_pt[37] | rom_instr_pt[64]
     | rom_instr_pt[65] | rom_instr_pt[69]
     | rom_instr_pt[126] | rom_instr_pt[130]
    );
assign count_src[0] =
    (rom_instr_pt[68] | rom_instr_pt[147]
     | rom_instr_pt[176] | rom_instr_pt[199]
    );
assign count_src[1] =
    (rom_instr_pt[68] | rom_instr_pt[176]
     | rom_instr_pt[196] | rom_instr_pt[199]
    );
assign count_src[2] =
    (rom_instr_pt[68] | rom_instr_pt[135]
     | rom_instr_pt[145] | rom_instr_pt[188]
     | rom_instr_pt[199]);
assign ext_rt =
    (rom_instr_pt[11] | rom_instr_pt[18]
     | rom_instr_pt[28] | rom_instr_pt[33]
     | rom_instr_pt[45] | rom_instr_pt[47]
     | rom_instr_pt[55] | rom_instr_pt[67]
     | rom_instr_pt[85] | rom_instr_pt[87]
     | rom_instr_pt[102] | rom_instr_pt[115]
     | rom_instr_pt[118] | rom_instr_pt[136]
     | rom_instr_pt[137] | rom_instr_pt[144]
     | rom_instr_pt[146] | rom_instr_pt[150]
     | rom_instr_pt[158] | rom_instr_pt[160]
     | rom_instr_pt[161] | rom_instr_pt[174]
     | rom_instr_pt[190] | rom_instr_pt[197]
    );
assign ext_s1 =
    (rom_instr_pt[33] | rom_instr_pt[36]
     | rom_instr_pt[45] | rom_instr_pt[55]
     | rom_instr_pt[63] | rom_instr_pt[67]
     | rom_instr_pt[74] | rom_instr_pt[85]
     | rom_instr_pt[96] | rom_instr_pt[101]
     | rom_instr_pt[115] | rom_instr_pt[118]
     | rom_instr_pt[135] | rom_instr_pt[136]
     | rom_instr_pt[137] | rom_instr_pt[144]
     | rom_instr_pt[150] | rom_instr_pt[151]
     | rom_instr_pt[152] | rom_instr_pt[157]
     | rom_instr_pt[160] | rom_instr_pt[173]
     | rom_instr_pt[179] | rom_instr_pt[182]
     | rom_instr_pt[185] | rom_instr_pt[189]
    );
assign ext_s2 =
    (rom_instr_pt[7] | rom_instr_pt[36]
     | rom_instr_pt[45] | rom_instr_pt[47]
     | rom_instr_pt[52] | rom_instr_pt[67]
     | rom_instr_pt[87] | rom_instr_pt[115]
     | rom_instr_pt[137] | rom_instr_pt[138]
     | rom_instr_pt[146] | rom_instr_pt[156]
     | rom_instr_pt[158] | rom_instr_pt[179]
     | rom_instr_pt[198]);
assign ext_s3 =
    (rom_instr_pt[22] | rom_instr_pt[116]
     | rom_instr_pt[161] | rom_instr_pt[168]
     | rom_instr_pt[182] | rom_instr_pt[193]
     | rom_instr_pt[197]);
assign sel0_5 =
    (rom_instr_pt[156]);
assign sel6_10[0] =
    (rom_instr_pt[97] | rom_instr_pt[120]
     | rom_instr_pt[122] | rom_instr_pt[128]
     | rom_instr_pt[159] | rom_instr_pt[162]
     | rom_instr_pt[175]);
assign sel6_10[1] =
    (rom_instr_pt[62] | rom_instr_pt[87]
     | rom_instr_pt[138] | rom_instr_pt[156]
     | rom_instr_pt[179] | rom_instr_pt[181]
     | rom_instr_pt[191]);
assign sel11_15[0] =
    (rom_instr_pt[36] | rom_instr_pt[63]
     | rom_instr_pt[101]);
assign sel11_15[1] =
    (rom_instr_pt[5] | rom_instr_pt[7]
     | rom_instr_pt[11] | rom_instr_pt[12]
     | rom_instr_pt[18] | rom_instr_pt[36]
     | rom_instr_pt[63] | rom_instr_pt[96]
     | rom_instr_pt[97] | rom_instr_pt[101]
     | rom_instr_pt[102] | rom_instr_pt[123]
     | rom_instr_pt[146] | rom_instr_pt[156]
     | rom_instr_pt[159] | rom_instr_pt[162]
     | rom_instr_pt[165] | rom_instr_pt[175]
    );
assign sel16_20[0] =
    (rom_instr_pt[174]);
assign sel16_20[1] =
    (rom_instr_pt[2] | rom_instr_pt[5]
     | rom_instr_pt[22] | rom_instr_pt[26]
     | rom_instr_pt[28] | rom_instr_pt[33]
     | rom_instr_pt[41] | rom_instr_pt[76]
     | rom_instr_pt[97] | rom_instr_pt[116]
     | rom_instr_pt[120] | rom_instr_pt[122]
     | rom_instr_pt[140] | rom_instr_pt[159]
     | rom_instr_pt[162] | rom_instr_pt[165]
     | rom_instr_pt[168] | rom_instr_pt[173]
     | rom_instr_pt[174] | rom_instr_pt[175]
    );
assign sel21_25[0] =
    1'b0;
assign sel21_25[1] =
    (rom_instr_pt[2] | rom_instr_pt[5]
     | rom_instr_pt[26] | rom_instr_pt[97]
     | rom_instr_pt[99] | rom_instr_pt[120]
     | rom_instr_pt[156] | rom_instr_pt[159]
     | rom_instr_pt[162] | rom_instr_pt[163]
     | rom_instr_pt[168]);
assign sel26_30 =
    (rom_instr_pt[2] | rom_instr_pt[5]
     | rom_instr_pt[26] | rom_instr_pt[97]
     | rom_instr_pt[99] | rom_instr_pt[120]
     | rom_instr_pt[156] | rom_instr_pt[159]
     | rom_instr_pt[162] | rom_instr_pt[163]
     | rom_instr_pt[168]);
assign sel31 =
    (rom_instr_pt[2] | rom_instr_pt[5]
     | rom_instr_pt[26] | rom_instr_pt[97]
     | rom_instr_pt[99] | rom_instr_pt[119]
     | rom_instr_pt[140] | rom_instr_pt[154]
     | rom_instr_pt[156] | rom_instr_pt[159]
     | rom_instr_pt[163]);
assign cr_bf2fxm =
    (rom_instr_pt[165]);
assign skip_cond =
    (rom_instr_pt[44] | rom_instr_pt[47]
     | rom_instr_pt[52] | rom_instr_pt[58]
     | rom_instr_pt[74] | rom_instr_pt[83]
     | rom_instr_pt[104] | rom_instr_pt[112]
     | rom_instr_pt[117] | rom_instr_pt[138]
    );
assign skip_zero =
    1'b0;
assign skip_nop =
    (rom_instr_pt[13] | rom_instr_pt[15]
     | rom_instr_pt[34] | rom_instr_pt[75]
     | rom_instr_pt[93] | rom_instr_pt[133]
     | rom_instr_pt[187]);
assign loop_addr[0] =
    (rom_instr_pt[200]);
assign loop_addr[1] =
    (rom_instr_pt[44] | rom_instr_pt[119]
     | rom_instr_pt[122] | rom_instr_pt[140]
     | rom_instr_pt[175] | rom_instr_pt[182]
     | rom_instr_pt[185] | rom_instr_pt[197]
    );
assign loop_addr[2] =
    (rom_instr_pt[36] | rom_instr_pt[45]
     | rom_instr_pt[58] | rom_instr_pt[67]
     | rom_instr_pt[75] | rom_instr_pt[115]
     | rom_instr_pt[119] | rom_instr_pt[122]
     | rom_instr_pt[133] | rom_instr_pt[140]
     | rom_instr_pt[157] | rom_instr_pt[185]
     | rom_instr_pt[187] | rom_instr_pt[189]
    );
assign loop_addr[3] =
    (rom_instr_pt[67] | rom_instr_pt[133]
     | rom_instr_pt[163] | rom_instr_pt[182]
     | rom_instr_pt[187] | rom_instr_pt[189]
     | rom_instr_pt[193] | rom_instr_pt[198]
    );
assign loop_addr[4] =
    (rom_instr_pt[75] | rom_instr_pt[115]
     | rom_instr_pt[133] | rom_instr_pt[140]
     | rom_instr_pt[151] | rom_instr_pt[157]
     | rom_instr_pt[197]);
assign loop_addr[5] =
    (rom_instr_pt[22] | rom_instr_pt[67]
     | rom_instr_pt[75] | rom_instr_pt[115]
     | rom_instr_pt[122] | rom_instr_pt[140]
     | rom_instr_pt[150] | rom_instr_pt[158]
     | rom_instr_pt[173] | rom_instr_pt[190]
     | rom_instr_pt[193]);
assign loop_addr[6] =
    (rom_instr_pt[67] | rom_instr_pt[115]
     | rom_instr_pt[119] | rom_instr_pt[122]
     | rom_instr_pt[140]);
assign loop_addr[7] =
    (rom_instr_pt[22] | rom_instr_pt[58]
     | rom_instr_pt[67] | rom_instr_pt[115]
     | rom_instr_pt[140] | rom_instr_pt[168]
     | rom_instr_pt[173] | rom_instr_pt[175]
     | rom_instr_pt[182]);
assign loop_addr[8] =
    (rom_instr_pt[22] | rom_instr_pt[45]
     | rom_instr_pt[58] | rom_instr_pt[67]
     | rom_instr_pt[75] | rom_instr_pt[133]
     | rom_instr_pt[140] | rom_instr_pt[157]
     | rom_instr_pt[158] | rom_instr_pt[163]
     | rom_instr_pt[168] | rom_instr_pt[173]
     | rom_instr_pt[182] | rom_instr_pt[193]
     | rom_instr_pt[198]);
assign loop_addr[9] =
    1'b0;
assign loop_init[0] =
    1'b0;
assign loop_init[1] =
    1'b0;
assign loop_init[2] =
    1'b0;
assign ep =
    (rom_instr_pt[7] | rom_instr_pt[22]
     | rom_instr_pt[41] | rom_instr_pt[116]
     | rom_instr_pt[146]);

//assign_end

   // Old FDIV/FSQRT
   //end generate;
   //| 1111000001    | 11111100001-----0000000000111100 0 - 0 - ---  1 0 1 1  0 00 10 00 00 0 0  0 0 - 0 ---------- --- -    | # fnmsub   s1,FB,s0,s0
   //| 1111000011    | 11111100011000010000100001111010 0 - 0 - ---  1 1 1 1  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # fmadd    s3,s1,s1,s1
   //| 1111000101    | 11111100000----------00010111100 0 - 0 - ---  1 0 0 1  0 00 10 11 00 0 0  0 0 - 0 ---------- --- -    | # fnmsub   s0,FB,s2,FA
   //| 1111000111    | 11111100000000010000000000110010 0 - 0 - ---  1 1 0 1  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # fmul     s0,s1,s0
   //| 1111001001    | 11111100011000000001000011111010 0 - 0 - ---  1 1 1 1  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # fmadd    s3,s0,s3,s2
   //| 1111001011    | 11111100010----------00011111100 0 - 0 - ---  1 0 0 1  0 00 10 11 00 0 0  0 0 - 0 ---------- --- -    | # fnmsub   s2,FB,s3,FA
   //| 1111001101    | 111111-----00001000000000010001- 1 - 0 - ---  0 1 1 1  0 01 00 00 00 0 1  0 0 - 0 ---------- --- -    | # fmul_uc  FT,s1,s0,s0  include s0 in 16-20
   //| 1111010001    | 11111100011-----0000000000111100 0 - 0 - ---  1 0 1 1  0 00 10 00 00 0 0  0 0 - 0 ---------- --- -    | # fnmsub   s3,FB,s0,s0
   //| 1111010011    | 11101100001000000000000011111010 0 - 0 - ---  1 1 1 1  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # fmadds   s1,s0,s3,s0
   //| 1111010101    | 11101100000----------00001111100 0 - 0 - ---  1 0 0 1  0 00 10 11 00 0 0  0 0 - 0 ---------- --- -    | # fnmsub   s0,FB,s1,FA
   //| 1111010111    | 11101100000----------00001111100 0 - 0 - ---  1 0 0 1  0 00 10 11 00 0 0  0 0 - 0 ---------- --- -    | # fnmsub   s0,FB,s1,FA
   //| 1111100001    | 11111100001000000000000000110010 0 - 0 - ---  1 1 0 1  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # fmul     s1,s0,s0,
   //| 1111100011    | 11111100000000010000100010111100 0 - 0 - ---  1 1 1 1  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # fnmsub   s0,s1,s2,s1
   //| 1111100101    | 11111100010000010000100000111010 0 - 0 - ---  1 1 1 1  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # fmadd    s2,s1,s0,s1
   //| 1111100111    | 11111100001000000001100010111010 0 - 0 - ---  1 1 1 1  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # fmadd    s1,s0,s2,s3
   //| 1111101001    | 1111110000000001-----00001111100 0 - 0 - ---  1 1 0 1  0 00 00 01 00 0 0  0 0 - 0 ---------- --- -    | # fnmsub   s0,s1,s1,FB
   //| 1111101011    | 1111110000000001-----00011111100 0 - 0 - ---  1 1 0 1  0 00 00 01 00 0 0  0 0 - 0 ---------- --- -    | # fnmsub   s0,s1,s3,FB
   //| 1111110001    | 11111100010000000000000000110010 0 - 0 - ---  1 1 0 1  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # fmul     s1,s0,s0,
   //| 1111110011    | 1111110000000011-----00011111100 0 - 0 - ---  1 1 0 1  0 00 00 01 00 0 0  0 0 - 0 ---------- --- -    | # fnmsub   s0,s2,s2,FB
   //| 1111110101    | 11101100011000000001100010111010 0 - 0 - ---  1 1 1 1  0 00 00 00 00 0 0  0 0 - 0 ---------- --- -    | # fmadds   s3,s0,s1,s2
   //| 1111110111    | 1110110001000011-----00011111100 0 - 0 - ---  1 1 0 1  0 00 00 01 00 0 0  0 0 - 0 ---------- --- -    | # fnmsubs  s2,s3,s3,FB
   //| 1111111001    | 111011-----00001000000000010001- 1 - 0 - ---  0 1 1 1  0 01 00 00 00 0 1  0 0 - 0 ---------- --- -    | # fmuls_uc FT,s1,s0,s0  include s0 in 16-20
   //32-bit core
   //c32: if (regmode = 5) generate begin
   //end generate;


   // ??? Do I want to optimize any terms?
   // ??? Which is better: on-off, or on-dc?
   // ??? Do we want to DC template fields not being used?

   assign rom_addr_d = rom_addr;

   assign rom_data = {template, ucode_end, ucode_end_early, loop_begin, loop_end, count_src, ext_rt, ext_s1, ext_s2, ext_s3, sel0_5, sel6_10, sel11_15, sel16_20, sel21_25, sel26_30, sel31, cr_bf2fxm, skip_cond, skip_zero, skip_nop, loop_addr, loop_init, ep};

   //---------------------------------------------------------------------
   // Latches
   //---------------------------------------------------------------------

   tri_rlmreg_p #(.WIDTH(10), .INIT(0), .NEEDS_SRESET(0)) rom_addr_latch(
      .vd(vdd),
      .gd(gnd),
      .nclk(nclk),
      .act(rom_act),
      .thold_b(pc_iu_func_sl_thold_0_b),
      .sg(pc_iu_sg_0),
      .force_t(force_t),
      .delay_lclkr(delay_lclkr),
      .mpw1_b(mpw1_b),
      .mpw2_b(mpw2_b),
      .d_mode(d_mode),
      .scin(siv[rom_addr_offset:rom_addr_offset + 10 - 1]),
      .scout(sov[rom_addr_offset:rom_addr_offset + 10 - 1]),
      .din(rom_addr_d),
      .dout(rom_addr_l2)
   );

   //---------------------------------------------------------------------
   // Scan
   //---------------------------------------------------------------------
   assign siv[0:scan_right] = {sov[1:scan_right], scan_in};
   assign scan_out = sov[0];

endmodule
