// © IBM Corp. 2020
// This softcore is licensed under and subject to the terms of the CC-BY 4.0
// license (https://creativecommons.org/licenses/by/4.0/legalcode). 
// Additional rights, including the right to physically implement a softcore 
// that is compliant with the required sections of the Power ISA 
// Specification, will be available at no cost via the OpenPOWER Foundation. 
// This README will be updated with additional information when OpenPOWER's 
// license is available.

// *!****************************************************************
// *! FILENAME    : tri_a2o.param
// *! DESCRIPTION : Constants for use throughout core
// *! CONTENTS    :
// *!
// *!****************************************************************

`ifndef _tri_vh_
`define _tri_vh_

`define  NCLK_WIDTH  6   // 0  1xClk, 1  Reset, 2  2xClk, 3  4xClk,  4  Even .5xClk,  5 Odd .5x Clk
//`define  EXPAND_TYPE  1

// Do NOT add any defines below this line
`endif  //_tri_vh_
